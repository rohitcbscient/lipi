b0VIM 8.0      ��`�t �  rohit                                   bhargav                                 ~rohit/my_git/lipi/adhyan/vla/20160409_analysis.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp"           j                            m       k                     G       �                     7                           ,       V                    C       �                    1       �                    4       �                    I       *                    :       s                    7       �                    1       �                    >                           >       S                    F       �                    =       �                    C                           8       W                    4       �                    ;       �                     ?       �             !       e       =                    &       �                           �             "       *       �             #                                  ?                           5       X                    B       �             	       @       �             
       ?                           @       N                    4       �                    ^       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     j       �  �  �  �  �  ~  U  ;    �  �  �  �  �  m  O  B  )    �  �  �  �  �  �  �  i  (    �  �  �  �  �  J  *  
  �  �  w  T  8     �
  �
  �
  G
  �	  �	  a	  R	  Q	  P	  +	  	  �  �  �  |  Z  =       �  �  �  n  L  *  �  �  �  �  \  @  (  �  �  �  O  �  �  i  Z  Y  X  =  *  �  �  �  �  c  G    �  �  �  �  i  E      �  �  �          def get_sunpy_maps(f):      return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data             maplist[i]=idl2sunpy_sdo(f[i],wave,inst)         if(inst=='AIA'):             maplist[i]=idl2sunpy_hmi(f[i])         if(inst=='HMI'):     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] def get_sunpy_maps_rot(f,wave,inst):      return sec     sec=ut.hms2sec_c(hhmmss)     hhmmss=' '+str(date.hour)+':'+str(date.minute)+':'+str(date.second)+'.'+str(date.microsecond/1.e6).split('.')[1]     date=mapp.date def produce_tstring(mapp):       return smp     smp = smap.Map(dat, header)     header['DSUN_OBS'] = sunpy.coordinates.get_sunearth_distance(header['DATE-OBS']).to(u.meter).value     header['RSUN_OBS'] = 958.11#sunpy.coordinates.sun.angular_radius(header['DATE-OBS']).value     header['RSUN_REF'] = sunpy.sun.constants.radius.value     header['HGLT_OBS'] = sunpy.coordinates.get_sun_B0(header['DATE-OBS']).value     header['HGLN_OBS'] = 0.     header['NAXIS2'], header['NAXIS1'] = dat.shape     header['NAXIS'] = 2     header['P_ANGLE'] = 0.0     header['waveunit'] = 'angstrom'     header['WAVELNTH'] = wave     header['INSTRUME'] = inst     header['TELESCOP'] = 'SDO'     header['CRPIX2'], header['CRPIX1'] = (np.array(dat.shape) + 1.0) / 2 + 0.5     header['CTYPE2'] = 'HPLT-TAN'     header['CTYPE1'] = 'HPLN-TAN'     header['CUNIT2'] = 'arcsec'     header['CUNIT1'] = 'arcsec'     header['DATE-OBS'] = Time(parser.parse(mp[5])).isot     header['CDELT2'] = mp[4]     header['CDELT1'] = mp[3]     header['CRVAL2'] = mp[2]     header['CRVAL1'] = mp[1]     header['EXPTIME'] = mp['dur']     header = {}     dat = np.nan_to_num(mp[0]) + 1e-6 # just to get rid of zeros     mp = mapstruc[keys[0]][0]     keys = list(mapstruc.keys())     mapstruc = readsav(mapsav) def idl2sunpy_sdo(mapsav,wave,inst):       return smp     smp = smap.Map(dat, header)     header['DSUN_OBS'] = sunpy.coordinates.get_sunearth_distance(header['DATE-OBS']).to(u.meter).value     header['RSUN_OBS'] = 958.11#sunpy.coordinates.sun.angular_radius(header['DATE-OBS']).value     header['RSUN_REF'] = sunpy.sun.constants.radius.value     header['HGLT_OBS'] = sunpy.coordinates.get_sun_B0(header['DATE-OBS']).value     header['HGLN_OBS'] = 0.     header['NAXIS2'], header['NAXIS1'] = dat.shape     header['NAXIS'] = 2     header['P_ANGLE'] = 0.0     header['TELESCOP'] = 'SDO/HMI'     header['CRPIX2'], header['CRPIX1'] = (np.array(dat.shape) + 1.0) / 2 + 0.5     header['CTYPE2'] = 'HPLT-TAN'     header['CTYPE1'] = 'HPLN-TAN'     header['CUNIT2'] = 'arcsec'     header['CUNIT1'] = 'arcsec'     header['DATE-OBS'] = Time(parser.parse(mp[5])).isot     header['CDELT2'] = mp[4]     header['CDELT1'] = mp[3]     header['CRVAL2'] = mp[2]     header['CRVAL1'] = mp[1]     header['EXPTIME'] = mp['dur']     header = {}     dat = np.nan_to_num(mp[0]) + 1e-6 # just to get rid of zeros     mp = mapstruc[keys[0]][0]     keys = list(mapstruc.keys())     mapstruc = readsav(mapsav) def idl2sunpy_hmi(mapsav):   import numpy as np from dateutil import parser from sunpy import sun import sunpy.map as smap import sunpy from astropy.time import Time from scipy.io import readsav import os import matplotlib.patches as patches from mpl_toolkits.axes_grid1 import make_axes_locatable import pickle import matplotlib as mpl from surya.utils import main as ut import astropy.units as u from astropy.coordinates import SkyCoord from sunpy.map import Map  from astropy.io import fits  import glob import sys import matplotlib.pyplot as plt import numpy as np ad  7   �     ^       �  �  �    t    �  �  p  -    �  �  �  �  p  8    �  �  b  "  �  �  B  �
  �
  x
  )
  �	  �	  p	  	  	  	  	  	  �  �  *            �  �  v  f  O  /       �  �  �  �  �  �  �  y  m  V  2      �  �  s  \  :  �  �  �  /    �  �  �  ~  s  r  c  Q  >  #    �  d  >  �  �  �  �  �                                                              plt.show()     ax2.set_ylabel('Amp')     ax2.plot(np.arange(150)/20.0,np.nanmean(ds_I2[10:20,:],axis=0),'o-')     ax1.set_ylabel('Frequency (GHz)')     ax2.set_xlabel('Time (s)')     ax1.imshow(np.log(ds_I2),aspect='auto',cmap='jet',extent=[time[0],7.5,freq[0],1.122],interpolation=None,origin=0,vmin=-3,vmax=1)     ax2=f.add_subplot(212)     ax1=f.add_subplot(211)     f=plt.figure() if(plot_full_ds): plot_full_ds=0  plt.show() ax2.set_xlabel('Time (HH:MM) UT') ax1.set_ylabel('Frequency (GHz)') ax2.set_xlim([0,600]) ax1.set_yticklabels([1.0,1.2,1.4,1.6,1.8,2.0]) ax1.set_yticks([0,100,200,300,400,500]) ax2.set_xticklabels(['18:40','18:41','18:42','18:43','18:44','18:45','18:46','18:47','18:48','18:49','18:50']) ax2.set_xticks([0,60,120,180,240,300,360,420,480,540,600]) ax2.plot(ds_feature2[10],'o-') ax1.imshow(ds_feature2,origin=0,vmin=0.01,vmax=0.8,aspect='auto') ax2=f.add_subplot(212,sharex=ax1) ax1=f.add_subplot(211) f=plt.figure()  #plt.imshow(np.log(ds_I1),aspect='auto',extent=[time[0],time[-1],freq[0],freq[-1]],cmap='jet',interpolation=None,origin=0,vmin=-3,vmax=1)  ds_feature2=ds_I[:,2585:2585+10*60] time_feature2=time[2585:2585+10*60] # 18:40:00 to 19:00:00 # Feature 2 #ds_I2=ds_I[:,2050:2200] #ds_I1=ds_I[:,:2680] # For feature 1  #   ds_I[:,i*120]=np.nan #for i in range(120): #ds_I=ds_I[:,771:] ds_I=0.5*(ds_LL+ds_RR) ds_RR=ds[1][0] ds_LL=ds[0][0] time=data['tim']-data['tim'][0] freq=data['freq']/1.e9 ds=data['spec'] data=np.load('sun_L_20160409.1s.ms.dspec.npz') plt.style.use('/home/i4ds1807205/scripts/general/plt_style.py') # Time from 17:59:56-22:57:52 sys.exit()   plt.show() compmap.plot() compmap.set_plot_settings(1,{'cmap':'gray','norm':mpl.colors.Normalize(vmin=-1.,vmax=1.),'origin':0}) compmap.set_levels(1,[10,20,30,40,50,60,70,80,90],percent=True) compmap=Map(map131[10],mapvla[0],composite=True)            plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs/aia1600_contour_'+str("%03d"%i)+'.png')     plt.title('VLA: '+v1.meta['date-obs'])     plt.text(401,50,'Contours: 15,18,21,27 MK',color='yellow')     plt.text(401,150,str(np.round(v3.meta['crval3']/1.e9,4))+' GHz',color='b')     plt.text(401,200,str(np.round(v2.meta['crval3']/1.e9,4))+' GHz',color='g')     plt.text(401,250,str(np.round(v1.meta['crval3']/1.e9,4))+' GHz',color='r')     plt.xlim([400,900]);plt.ylim([50,550])     v3.draw_contours(levels=lev3,colors='b',linewidths=3,extent=p.get_extent())     v2.draw_contours(levels=lev2,colors='g',linewidths=3,extent=p.get_extent())     v1.draw_contours(levels=lev1,colors='r',linewidths=3,extent=p.get_extent())     lev3=(3.e7/v3.data.max())*np.array([50,60,70,90])*u.percent     lev2=(3.e7/v2.data.max())*np.array([50,60,70,90])*u.percent     lev1=(3.e7/v1.data.max())*np.array([50,60,70,90])*u.percent     v3=allmaps['vla']['mapvla'][119*freq_id[2]+i]     v2=allmaps['vla']['mapvla'][119*freq_id[1]+i]     v1=allmaps['vla']['mapvla'][119*freq_id[0]+i]     p=allmaps['aia1600']['map1600'][tidx1600[i]].plot() for i in range(119):      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia131_contour_'+str("%03d"%i)+'.png')     plt.show()     #plt.xlim([400,900]);plt.ylim([50,550])     plt.text(401,50,'Contours: 1.5,1.8,2.1,2.7 MK',color='yellow')     plt.text(401,250,str(np.round(v1.meta['crval3']/1.e9,4))+' GHz',color='r')     compmap.plot()     compmap.set_levels(1,[30,40,50,60,70,80,90],percent=True)     compmap=Map(allmaps['aia171']['map171'][tidx171[i]],allmaps['vla']['mapvla'][i],composite=True)     i=1400 for i in range(1):      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia1600_contour_'+str("%03d"%i)+'.png') ad  p
  �
            �  �  �  �  �  i  +    0  �  s  ;  �  �  m  b  a  `  B  )    �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      dd=v;dd.data[np.isnan(dd.data)]=0 cc=allmaps['aia171']['map171'][10] ax0 = f.add_subplot(111) f=plt.figure(figsize=(10,10))   plt.show() ax0.set_xlim([-900,-700]),ax0.set_ylim([100,300]) #ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow') #ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r') ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia]) ax0.set_title('AIA 171 $\AA$:18:42:10 UT VLA: 18:44:43.00-18:44:43.05 UT') dd.draw_contours(levels=lev1,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2) lev1=np.array([60,70,80,90])*u.percent #lev1=(1.5e7/dd.data.max())*np.array([60,70,80,90])*u.percent p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2) dd=v;dd.data[np.isnan(dd.data)]=0 cc=allmaps['aia171']['map171'][10] ax0 = f.add_subplot(111) f=plt.figure(figsize=(10,10)) ad  ?  �     &       �  b  :  �  �  x  2  �  I  �  w    �  �  -    �
  F
  �	  �	  �	  �	  s	  d	  	  �  �  n  G  �  w  T  I  H  �    �  �    �  �     �    X  �    �  �  C  �  �  �  �  �  �  }  Z  8                                                      dd=v;dd.data[np.isnan(dd.data)]=0 cc=allmaps['aia171']['map171'][10] ax0 = f.add_subplot(111) f=plt.figure(figsize=(10,10))   plt.show() ax0.set_xlim([-900,-700]),ax0.set_ylim([100,300]) #ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow') #ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r') ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia]) ax0.set_title('AIA 171 $\AA$:18:42:10 UT VLA: 18:44:43.00-18:44:43.05 UT') dd.draw_contours(levels=lev1,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2) lev1=np.array([60,70,80,90])*u.percent #lev1=(1.5e7/dd.data.max())*np.array([60,70,80,90])*u.percent p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aslistvla_rr=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_6/*spw.6_16-31*FITS'));v6=Map(listvla_rr[860]);v6.data[np.isnan(v6.data)]=0 listvla_rr=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_4/*spw.4_16-31*FITS'));v4=Map(listvla_rr[860]);v4.data[np.isnan(v4.data)]=0 listvla_rr=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_2/*spw.2_16-31*FITS'));v2=Map(listvla_rr[860]);v2.data[np.isnan(v2.data)]=0 listvla_rr=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_0/*spw.0_16-31*FITS'));v=Map(listvla_rr[860]);v.data[np.isnan(v.data)]=0  plt.show() ax.legend(loc=4);ax1.legend(loc=2) ax.set_ylabel('Flux (W/m$^2$)');ax1.set_ylabel('Flux (W/m$^2$)');ax.set_xlabel('Time (HH:MM UT)') ax.set_xticklabels(['18:30','18:33','18:36','18:39','18:42','18:45','18:48','18:51','18:54','18:57','19:00']) ax.set_xticks(np.arange(11)*180+66601) ax.axvline(x=67798,linestyle='--',color='k') ax.axvline(x=67200,linestyle='--',color='k') #ax.plot(gtime[292:585]-600+67200,gf0540[292:585],'o-',color='g',label='0.5-4.0$\AA$') ax1.plot(gtime-600+67200,gf1080,'o-',color='b',label='1.0-8.0$\AA$') ax1=ax.twinx() ax.plot(gtime-600+67200,gf0540,'o-',color='g',label='0.5-4.0$\AA$') f,ax=plt.subplots(1,1)      plt.show()     ax[2].set_xlim([67200.,67560.]);ax[2].set_ylabel('Flux (W/m$^2$)');ax2.set_ylabel('Flux (W/m$^2$)')     ax[1].set_ylabel('Amplitude');ax[2].set_xlabel('Time (HH:MM UT)')#;ax1.set_ylabel('')     ax2.plot(gtime[292:585]-600+67200,gf1080[292:585],'o-',label='1.0-8.0$\AA$');ax[2].legend(loc=4);ax2.legend(loc=2)     ax2=ax[2].twinx()     ax[2].plot(gtime[292:585]-600+67200,gf0540[292:585],'o-',color='g',label='0.5-4.0$\AA$')     ax[1].legend(loc=2,prop={'size':15})     #plt.ylabel('T$_{B}$ ($\\times10^{5}$ (K))');plt.xlabel('Time (HH:MM UT)')     ax[1].set_xticklabels(['18:40','18:41','18:42','18:43','18:44','18:45','18:46','18:47','18:48','18:49','18:50'])     ax[1].set_xticks(np.arange(11)*60+67212-11)     #ax1.plot(np.hstack((np.array(qstimevla)[:,0],np.array(timevla_all)[0:2000])),np.hstack((np.array(qsTbr_r1),Tbr_r1[1]))/1.e8,'-',color='k',label='1.077 GHz')     ax[1].plot(fmtime[14244:14332],fmrate[14244:14332:,0:20].mean(axis=1)/200,'o-',color='orange',label='FERMI')     ax[1].plot(qstimevla[0][0]+np.arange(7200)*0.05,ds_LL1[0:128].mean(axis=0)/120,'-',color='k',label='0.99-1.25 GHz')     ax[1].plot(time1600,ts1600-ts1600[1],'o-',label='AIA 1600 $\AA$')     ax[1].plot(time335,ts335-ts335[1],'o-',label='AIA 335 $\AA$')     ax[1].plot(time131,ts131-ts131[1],'o-',label='AIA 131 $\AA$')     ax[1].plot(time94,ts94-ts94[1],'o-',label='AIA 94 $\AA$')     ax[0].set_ylabel('Frequency (GHz)')     ax[0].imshow(ds_LL1,aspect='auto',origin=0,cmap='YlGnBu',vmin=10,vmax=80,extent=[67200.0,67560.,freq[0],freq[-1]])     f,ax=plt.subplots(3,1,sharex=True) ad     #     ?       �  y  x  d  M  $  �  �  p  =  �  �  X    �  �  V  +  �  �  �  y  P    �
  j
  .
  �	  �	  ,	  	  	  	  �  �  �  y  O  o  -  �  �  �  �  �  L  +    #  �  �  �  \  |  :     �  �  �  �  m  I  #  "                     f=plt.figure(figsize=(10,10))     for i in range(1,len(maphmir)): if(plot_base_hmi_movie): plot_run_hmi_movie=1          plt.close()         plt.savefig('/media/rohit/VLA/20160409/pngs/aia_'+str("%03d"%i)+'.png')         ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmaps['aia335']['map335'][i]         ax0 = f.add_subplot(224)         ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmaps['aia94']['map94'][i]         ax0 = f.add_subplot(223)         ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmaps['aia171']['map171'][i]         ax0 = f.add_subplot(222)         ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmaps['aia131']['map131'][i]         ax0 = f.add_subplot(221)         f=plt.figure(figsize=(10,10))     for i in range(len(allmaps['aia131']['data131'])): if(plot_aia_movie): plot_aia_movie=1      plt.show()     #ax[1].set_xticks([0,10,20,30]);ax[1].set_xticklabels([freq[0],freq[10],freq[20],freq[30]])     ax[1].legend();ax[1].set_ylabel('Source size (arcsec$^{2}$)');ax[1].set_xlabel('Frequency (GHz)')     ax[1].plot(freq,Tb_mean_r1[:,51],'o-',label='18:44:51')     ax[1].plot(freq,Tb_mean_r1[:,46],'o-',label='18:44:46')     ax[0].legend();ax[0].set_ylabel('Source size (arcsec$^{2}$)');ax[0].set_xlabel('Frequency (GHz)')     ax[0].plot(freq,vlasize_fwhm[0,:,51],'o-',label='18:44:51')     ax[0].plot(freq,vlasize_fwhm[0,:,46],'o-',label='18:44:46')     fig,ax=plt.subplots(2,1,sharex=True) if(plot_vlasize_freq): plot_vlasize_freq=1     plt.show()     ax[0].set_ylabel('Frequency (GHz)');ax[1].set_ylabel('T$_{B}$ (MK)');ax[2].set_ylabel('Source size (arcsec$^{2}$)')     ax[2].set_xlabel('Time (HH:MM:SS UT)')     ax[2].set_xticks([0,30,60,90,120]);ax[2].set_xticklabels(['18:44:00','18:44:30','18:45:00','18:45:30','18:46:00'])     ax[2].legend()     ax[2].plot(vlasize_fwhm[3,10],'o',label='90% Contours')     ax[2].plot(vlasize_fwhm[2,10],'o',label='70% Contours')     ax[2].plot(vlasize_fwhm[0,10],'o',label='50% Contours')     ax[1].plot(Tb_mean_r1[10]/1.e6,'o-',label='1.077 GHz');ax[1].legend()     ax[0].set_yticks([0,10,20,30]);ax[0].set_yticklabels([freq[0],freq[10],freq[20],freq[30]])     fig.colorbar(im0,cax=cax,label='T$_{B}$ (MK)')     cax = divider.append_axes('right', size='5%', pad=0.05)     divider = make_axes_locatable(ax[0])     im0=ax[0].imshow(Tb_mean_r1/1.e6,origin=0,cmap='jet',interpolation='None')     fig,ax=plt.subplots(3,1,sharex=True) if(plot_vlasize_fwhm): plot_vlasize_fwhm=1      plt.show()     ax[0].set_ylabel('Frequency (GHz)');ax[1].set_ylabel('T$_{B}$ (MK)');ax[2].set_ylabel('Source size (arcsec$^{2}$)') ad          5       �  �  �  �  !  �  �  ~  }  g  N  ,    �  �  �  �  %  �
  �
  �
  �
  o
  Z
   
  �	  �	  �	  �  i    �  �  �  n    �  �  �  w    �  �  �  ~    �  �  �  �  z  A                                             p=allmaps['aia1600']['map1600'][i].plot()     for i in range(len(allmaps['aia1600']['data1600'])): if(plot_euv1600_movie): plot_euv1600_movie=1          plt.close()         plt.savefig('/media/rohit/VLA/20160409/pngs/base_zoom_aia_'+str("%03d"%i)+'.png')         ax0.set_xlim([-800,-730]);ax0.set_ylim([200,270]);ax0.plot([-778,-778],[245,268],'o',color='k')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-10,vmax=10,cmap='coolwarm')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmapsb['aiab335']['mapb335'][i]         ax0 = f.add_subplot(224)         ax0.set_xlim([-800,-730]);ax0.set_ylim([200,270]);ax0.plot([-778,-778],[245,268],'o',color='k')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-10,vmax=10,cmap='coolwarm')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmapsb['aiab94']['mapb94'][i]         ax0 = f.add_subplot(223)         ax0.set_xlim([-800,-730]);ax0.set_ylim([200,270]);ax0.plot([-778,-778],[245,268],'o',color='k')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-150,vmax=150,cmap='coolwarm')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmapsb['aiab171']['mapb171'][i]         ax0 = f.add_subplot(222)         ax0.set_xlim([-800,-730]);ax0.set_ylim([200,270]);ax0.plot([-778,-778],[245,268],'o',color='k')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-20,vmax=20,cmap='coolwarm')         xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)         cc=allmapsb['aiab131']['mapb131'][i]         ax0 = f.add_subplot(221)         f=plt.figure(figsize=(10,10))     for i in range(len(allmapsb['aiab171']['datab171'])): if(plot_base_movie): plot_base_movie=1          plt.close()         plt.savefig('/media/rohit/VLA/20160409/pngs/hmib1_'+str("%03d"%i)+'.png')         f.colorbar(p,orientation='horizontal',label='B (G)')         ax0.set_xlim([-800,-730]);ax0.set_ylim([200,270]);ax0.plot([-778,-778],[245,268],'o',color='cyan')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-150,vmax=150,cmap='binary')         xlaia=cc.center.Tx.value-0.5*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.5*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.5*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.5*int(cc.data.shape[0]/2)         cc=maphmib[i]         ax0 = f.add_subplot(111)         f=plt.figure(figsize=(10,10))     for i in range(len(maphmib)): if(plot_base_hmi_movie): plot_base_hmi_movie=1          plt.close()         plt.savefig('/media/rohit/VLA/20160409/pngs/hmir2_'+str("%03d"%i)+'.png')         f.colorbar(p,orientation='horizontal',label='B (G)')         ax0.set_xlim([-800,-730]);ax0.set_ylim([230,300]);ax0.plot([-778,-778],[245,268],'o',color='cyan')         p=cc.plot(extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-80,vmax=80,cmap='binary')         xlaia=cc.center.Tx.value-0.5*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.5*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.5*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.5*int(cc.data.shape[0]/2)         cc=maphmir[i]         ax0 = f.add_subplot(111) ad     7     B       �  }  i  h  g  U  B  7     �  �  x  D    �  �  V    �  d  8  �  �  I    �
  �
  p
  `
  _
  �	  l	  �  y  x  t  ^  <    �  �  �  �  @    0  �  b  &  �  �  *    �  �  V  �  �  �  �  �  �  �  �  r  7  6                         ax0.plot(x,ycimax[i],'o',color='red',label='Stokes I')     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(20, 10))     x=np.arange(2000)*0.05 for i in range(32): i=0       plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia131_contour_Tb_'+str("%03d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('Median Amplitude')     ax1.axvline(x=i*0.05,color='k')     ax1.plot(np.arange(2400)*0.05,ds[0].mean(axis=0)[0],'-',label='1.077 GHz')     ax1 = f.add_subplot(212)     #ax0.text(-1200,50,'Contours: 20%, 30%, 40%, 50%, 60%, 70%, 80%, 90%',color='yellow')     ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow')     ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r')     ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd.draw_contours(levels=lev1,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2)     #lev1=np.array([20,30,40,50,60,70,80,90])*u.percent     lev1=(1.5e7/dd.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     dd=allmaps['vla']['mapvla'][i];dd.data[np.isnan(dd.data)]=0     cc=allmaps['aia131']['map131'][tidx131[i]]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(6, 10)) for i in range(2399): i=0  #xrpix=cc.world_to_pixel(yr).x.value;yrpix=cc.world_to_pixel(yr).y.value #yr = SkyCoord(dd.center.Tx.value+0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value+0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec)) #xlpix=cc.world_to_pixel(xl).x.value;ylpix=cc.world_to_pixel(xl).y.value #xl = SkyCoord(dd.center.Tx.value-0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value-0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec))      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia131_contour_'+str("%03d"%i)+'.png')     plt.show()     plt.title('VLA: '+v1.meta['date-obs'])     plt.text(401,50,'Contours: 1.5,1.8,2.1,2.7 MK',color='yellow')     #plt.text(401,150,str(np.round(v3.meta['crval3']/1.e9,4))+' GHz',color='b')     #plt.text(401,200,str(np.round(v2.meta['crval3']/1.e9,4))+' GHz',color='g')     plt.text(401,250,str(np.round(v1.meta['crval3']/1.e9,4))+' GHz',color='r')     #plt.xlim([400,900]);plt.ylim([50,550])     #v3.draw_contours(levels=lev3,colors='b',linewidths=3,extent=p.get_extent())     #v2.draw_contours(levels=lev2,colors='g',linewidths=3,extent=p.get_extent())     v1.draw_contours(levels=lev1,colors='r',linewidths=3,extent=p.get_extent())     #lev3=(3.e7/v3.data.max())*np.array([50,60,70,90])*u.percent     #lev2=(3.e7/v2.data.max())*np.array([50,60,70,90])*u.percent     lev1=np.array([50,60,70,90])*u.percent     #lev1=(1.e7/v1.data.max())*np.array([50,60,70,90])*u.percent     #v3=allmaps['vla']['mapvla'][2399*freq_id[2]+i]     #v2=allmaps['vla']['mapvla'][2399*freq_id[1]+i]     v1.data[np.isnan(v1.data)]=0     v1=allmaps['vla']['mapvla'][2399*freq_id[0]+i]     p=allmaps['aia1600']['map1600'][tidx131[i]].plot()     i=1400 for i in range(1): freq_id=[0,15,30]           plt.close()         plt.savefig('/media/rohit/VLA/20160409/pngs/aia1600_'+str("%03d"%i)+'.png')         plt.xlim([400,900]);plt.ylim([50,550]) ad  =   Y     @       �  �      �  �  '  �  �  �  �  �  �  �  q  M  *    �  �  {  D  h  !  S
  �	  .	  �  �  �  S  6  �  �  f  3     �  �  �  B  �  �  �  �  �  �  �  P  �  �  �  �  �  ^    �  �  r  #  �  �  �  Y  X                                                                   ax1.set_xlabel('Time (sec)');ax1.set_ylabel('$T_B$ (MK)')     ax1.axvline(x=x[50],color='k');ax1.set_ylim(0,100)     ax1.legend(loc=2)     ax1.plot(x[50],y[i+50]/1.e6,'o',color='red',markersize=10)     ax1.plot(x,y[i:i+100]/1.e6,'o-',markersize=5,label='Region 1 (0.994 GHz)')     ax1 = f.add_subplot(212)     ax0.set_xlim([-810,-750]);ax0.set_ylim([220,280])     #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     ax0.plot(centx[i+40:i+50],centy[i+40:i+50],'o',color='red')     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     ax0 = f.add_subplot(211)     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     cc=allmaps['aia171']['map171'][tidx171[i]]     f=plt.figure(figsize=(10, 15))     centx=np.hstack((np.array(qsxcr90),xcr90[1]));centy=np.hstack((np.array(qsycr90),ycr90[1]))     y=np.hstack((np.array(qsTbr_r1),Tbr_r1[1]))     x=np.arange(6799)[i:i+100]*0.05 for i in range(2399,6799): i=0      plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms_spw0/centroid_llrr_'+str("%04d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('$T_B$ (MK)')     ax1.axvline(x=x[50],color='k');ax1.set_ylim(0,100)     ax1.legend(loc=2)     #ax1.plot(x,Tb_r[4]/1.e6,'-',label='Region 5')     #ax1.plot(x,Tb_r[3]/1.e6,'-',label='Region 4')     #ax1.plot(x,Tb_r[2]/1.e6,'-',label='Region 3')     #ax1.plot(x,Tb_r[1]/1.e6,'-',label='Region 2')     ax1.plot(x[50],TbRRr1[i+50][0]/1.e6,'o',color='red',markersize=10)     ax1.plot(x,TbRRr1[i:i+100,0]/1.e6,'o-',markersize=5,label='Region 1 (0.994 GHz)')     ax1 = f.add_subplot(212)     f.colorbar(im0,label='(RR) Frequency (GHz)')     ax0.set_xlim([-810,-750]);ax0.set_ylim([220,280])     #ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])     #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     im0=ax0.scatter(xcr90[i+50].reshape(1,32).mean(axis=0)[0:16],ycr90[i+50].reshape(1,32).mean(axis=0)[0:16],c=freq.reshape(1,32).mean(axis=0)[0:16],s=40,cmap=plt.cm.get_cmap('spring'),edgecolors='none')     #im0=ax0.scatter(xcl90[i+50].reshape(1,32).mean(axis=0)[0:16],ycl90[i+50].reshape(1,32).mean(axis=0)[0:16],c=freq.reshape(1,32).mean(axis=0)[0:16],s=40,cmap=plt.cm.get_cmap('winter'),edgecolors='none')     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     #dd=mapvla_v[i+50][0];dd.data[np.isnan(dd.data)]=0     #cc=allmaps['aia171']['map171'][tidx171[i]]     cc=allmaps['aia171']['map171'][tidx171[i]]     #cc=allmapsb['aiab171']['mapb171'][tidx171[i]]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(10, 15))     x=np.arange(2000)[i:i+100]*0.05 for i in range(1900): i=0  ################ Plot centroids on AIA      plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/spec_max/stokes_I_'+str("%04d"%i)+'.png')     ax2=ax1.twinx();ax2.plot(x,maxTbi[i]/1.e6,'-',color='black');ax2.set_ylabel('T$_B$ (MK)')     ax0.axhline(y=255,linestyle='--',color='black')     ax1.set_ylim(-30,30);ax0.set_ylim(235,275);ax0.legend();ax0.set_title(str(freq[i])+' GHz')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('Solar-Y (arcsec)');ax0.set_ylabel('Solar-Y (arcsec)')     ax1.plot(x,ycimax[i]-ycvmax[i],'o')     ax1 = f.add_subplot(212)     ax0.plot(x,ycvmax[i],'o',color='blue',label='Stokes V') ad     2     ?       �  �    ~  }  ^  ;  c  J    �  E  �  �  �  �  �  �  �  �  _  <    �  �  �  V  z
  3
  8	  6  �  �  j  4    �  z  G    �  �  �  a  #  �  �  �  �  �  �  e  B  %  �  �  �  ]  �  :  �  o  2  1                                #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     im0=ax0.scatter(xcvmax[:25,i],ycvmax[:25,i],c=freq[:25],s=40,cmap=plt.cm.get_cmap('RdYlBu'),edgecolors='none')     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     dd=mapvla_v[i+50][0];dd.data[np.isnan(dd.data)]=0     #cc=allmaps['aia171']['map171'][tidx171[i]]     cc=allmaps['aia171']['map171'][tidx171[i]]     #cc=allmapsb['aiab171']['mapb171'][tidx171[i]]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(10, 15))     x=np.arange(2000)[i:i+100]*0.05 for i in range(1900): i=0      plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms_spw0/centroid_llrr1_'+str("%04d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('$T_B$ (MK)')     ax1.axvline(x=x[50],color='k');ax1.set_ylim(0,100)     ax1.legend(loc=2)     #ax1.plot(x,Tb_r[4]/1.e6,'-',label='Region 5')     #ax1.plot(x,Tb_r[3]/1.e6,'-',label='Region 4')     #ax1.plot(x,Tb_r[2]/1.e6,'-',label='Region 3')     #ax1.plot(x,Tb_r[1]/1.e6,'-',label='Region 2')     ax1.plot(x[50],TbRRr1[i+50][0]/1.e6,'o',color='red',markersize=10)     ax1.plot(x,TbRRr1[i:i+100,0]/1.e6,'o-',markersize=5,label='Region 1 (0.994 GHz)')     ax1 = f.add_subplot(212)     ax0.set_xlim([-810,-750]);ax0.set_ylim([220,280])     #ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])     #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     im0=ax0.errorbar(xcRR90[i+50].reshape(1,32).mean(axis=0)[0:16].mean(),ycRR90[i+50].reshape(1,32).mean(axis=0)[0:16].mean(),xerr=xcRR90[i+50].reshape(1,32).mean(axis=0)[0:16].std(),yerr=ycRR90[i+50].reshape(1,32).mean(axis=0)[0:16].std(),color='magenta')     im0=ax0.errorbar(xcLL90[i+50].reshape(1,32).mean(axis=0)[0:6].mean(),ycLL90[i+50].reshape(1,32).mean(axis=0)[0:6].mean(),xerr=xcLL90[i+50].reshape(1,32).mean(axis=0)[0:6].std(),yerr=ycLL90[i+50].reshape(1,32).mean(axis=0)[0:6].std(),color='blue')     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     #dd=mapvla_v[i+50][0];dd.data[np.isnan(dd.data)]=0     #cc=allmaps['aia171']['map171'][tidx171[i]]     cc=allmaps['aia171']['map171'][tidx171[i]]     #cc=allmapsb['aiab171']['mapb171'][tidx171[i]]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(10, 15))     x=np.arange(2000)[i:i+100]*0.05 for i in range(1900): i=0   plt.show() ax0.set_xlim([-810,-750]);ax0.set_ylim([220,280]) ax0.legend() ax0.plot(centx[5000:],centy[5000:],'o',color='r',alpha=0.2,label='18:48:10 to 18:49:40 UT') ax0.plot(centx[2000:5000],centy[2000:5000],'o',color='g',alpha=0.2,label='18:45:40 to 18:48:10 UT') ax0.plot(centx[0:2000],centy[0:2000],'o',color='b',alpha=0.2,label='18:44:00 to 18:45:40 UT') p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') ax0 = f.add_subplot(111) xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2) cc=allmaps['aia171']['map171'][10] f=plt.figure(figsize=(15, 15))       plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms_spw0_qs/centroid_llrr_'+str("%04d"%i)+'.png') ad     0     @       �  �  g  J  �  �  }  J    �  �  �  Z  �  �  �  �  �  �  �  �  c  0    �  �  �
  x
  
  �	  �	  �  <  �  �  p  :  �  �  ?  �  �  &  �  ]  �  �  �  I    �  �  }  g  1  �  �  ~  n  m  l  h  R  0  /                          f=plt.figure(figsize=(6, 10)) for i in range(2399): i=0       plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms_spw0/regions_contour_base_'+str("%04d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('$T_B$ (MK)')     ax1.axvline(x=x[50],color='k');ax1.set_ylim(0,50)     ax1.legend(loc=2)     #ax1.plot(x,Tb_r[4]/1.e6,'-',label='Region 5')     #ax1.plot(x,Tb_r[3]/1.e6,'-',label='Region 4')     #ax1.plot(x,Tb_r[2]/1.e6,'-',label='Region 3')     #ax1.plot(x,Tb_r[1]/1.e6,'-',label='Region 2')     ax1.plot(x[50],Tb_r[0][i+50]/1.e6,'o',color='red',markersize=10)     ax1.plot(x,Tb_r[0][i:i+100]/1.e6,'o-',markersize=5,label='Region 1')     ax1 = f.add_subplot(212)     #ax0.add_patch(patches.Rectangle((-831,175),40,40,linewidth=5,edgecolor='magenta',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-961,195),40,40,linewidth=5,edgecolor='cyan',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-881,175),40,40,linewidth=5,edgecolor='r',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-841,265),20,20,linewidth=5,edgecolor='g',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-781,233),40,40,linewidth=5,edgecolor='b',facecolor='none'))     #ax0.text(-990,64,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow')     #ax0.text(-990,64,'Contours: 20%, 30%, 40%,50%, 60%, 70%, 80%, 90%',color='yellow')     #ax0.text(-1200,50,'Contours: 0.6,0.75,0.9,1.0,1.2,1.3 MK',color='yellow')     ax0.text(-830,210,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='white')     ax0.set_xlim([-830,-730]);ax0.set_ylim([200,300])     #ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350])     #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd.draw_contours(levels=lev1,colors='black',linewidths=1,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2)     lev1=np.array([50,60,70,80,90,99])*u.percent     #lev1=(1.5e7/dd.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent     #p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-150,vmax=150,cmap='coolwarm')     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     dd=mapvla_v[i+50][0];dd.data[np.isnan(dd.data)]=0     #cc=allmaps['aia171']['map171'][tidx171[i]]     cc=allmaps['aia171']['map171'][tidx171[i]]     #cc=allmapsb['aiab171']['mapb171'][tidx171[i]]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(6, 10))     x=np.arange(2000)[i:i+100]*0.05 for i in range(1900): i=0      plt.close()     f.clear()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms_spw0/centroid_'+str("%04d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('$T_B$ (MK)')     ax1.axvline(x=x[50],color='k');ax1.set_ylim(0,50)     ax1.legend(loc=2)     #ax1.plot(x,Tb_r[4]/1.e6,'-',label='Region 5')     #ax1.plot(x,Tb_r[3]/1.e6,'-',label='Region 4')     #ax1.plot(x,Tb_r[2]/1.e6,'-',label='Region 3')     #ax1.plot(x,Tb_r[1]/1.e6,'-',label='Region 2')     ax1.plot(x[50],Tb_r[0][i+50]/1.e6,'o',color='red',markersize=10)     ax1.plot(x,Tb_r[0][i:i+100]/1.e6,'o-',markersize=5,label='Region 1 (0.994 GHz)')     ax1 = f.add_subplot(212)     f.colorbar(im0,label='Frequency (GHz)')     ax0.set_xlim([-830,-730]);ax0.set_ylim([200,300])     #ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,350]) ad  5   !     4       �  �  t  �  Q    �    �  8  �  �  ^    �
  �
  �
  @
  �	  �	  �	  �	  �	  L	  <	  �  H  �  O    �  Y    �  �  /        �  �  �  C  �  J  �  Q  �  �  [  0  !                                                              plt.show()     plt.xlim([400,900]);plt.ylim([50,550])     plt.text(401,50,'Contours: 0.6,0.75,0.9,1.0,1.2,1.3 MK',color='yellow')     plt.text(401,250,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r')     dd.draw_contours(levels=lev1,colors='r',linewidths=3,extent=[xlpix,xrpix,ylpix,yrpix])     xrpix=cc.world_to_pixel(yr).x.value;yrpix=cc.world_to_pixel(yr).y.value     yr = SkyCoord(dd.center.Tx.value+0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value+0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec))     xlpix=cc.world_to_pixel(xl).x.value;ylpix=cc.world_to_pixel(xl).y.value     xl = SkyCoord(dd.center.Tx.value-0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value-0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec))     lev1=(1.5e7/dd.data.max())*np.array([40,50,60,70,80,90])*u.percent     p=cc.plot()     dd=allmaps['vla']['mapvla'][i];dd.data[np.isnan(dd.data)]=0     cc=allmaps['aia1600']['map1600'][tidx131[i]] for i in range(1):      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia1600_contour_'+str("%03d"%i)+'.png')     plt.xlim([400,900]);plt.ylim([50,550])     plt.title('AIA 1600 $\AA$:'+timstr_1600[tidx131[i]]+' VLA: '+timstr_vla[i]+' UT')     plt.text(401,50,'Contours: 0.6,0.75,0.9,1.0,1.2,1.3 MK',color='yellow')     plt.text(401,250,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r')     dd.draw_contours(levels=lev1,colors='r',linewidths=3,extent=[xlpix,xrpix,ylpix,yrpix])     xrpix=cc.world_to_pixel(yr).x.value;yrpix=cc.world_to_pixel(yr).y.value     yr = SkyCoord(dd.center.Tx.value+0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value+0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec))     xlpix=cc.world_to_pixel(xl).x.value;ylpix=cc.world_to_pixel(xl).y.value     xl = SkyCoord(dd.center.Tx.value-0.5*(2.0/0.6)*dd.data.shape[0],dd.center.Ty.value-0.5*(2.0/0.6)*dd.data.shape[1], frame=cc.coordinate_frame, unit=(u.arcsec, u.arcsec))     lev1=(1.5e7/dd.data.max())*np.array([40,50,60,70,80,90])*u.percent     p=cc.plot()     dd=allmaps['vla']['mapvla'][i];dd.data[np.isnan(dd.data)]=0     cc=allmaps['aia1600']['map1600'][tidx131[i]] for i in range(2399):      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_50ms/aia171_contour_'+str("%03d"%i)+'.png')     ax1.set_xlabel('Time (sec)');ax1.set_ylabel('Median Amplitude')     ax1.axvline(x=i*0.05,color='k')     ax1.plot(np.arange(2400)*0.05,ds[0].mean(axis=0)[0],'-',label='1.077 GHz')     ax1 = f.add_subplot(212)     ax0.text(-1200,50,'Contours: 50%, 60%, 70%, 80%, 90%',color='yellow')     #ax0.text(-1200,50,'Contours: 0.6,0.75,0.9,1.0,1.2,1.3 MK',color='yellow')     ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r')     ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd.draw_contours(levels=lev1,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2)     lev1=np.array([50,60,70,80,90])*u.percent     #lev1=(1.5e7/dd.data.max())*np.array([50,60,70,80,90])*u.percent     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     dd=allmaps['vla']['mapvla'][i];dd.data[np.isnan(dd.data)]=0     cc=allmaps['aia171']['map171'][tidx131[i]]     ax0 = f.add_subplot(211) ad  A        m       �  �  �  {  W  +    �  �  �  �  v  _  F    �  �  �  �  q  S  .      �  �  �  m  Q  -    �  �  �  �  �  �  J  1    �
  �
  y
  >
  
  �	  �	  �	  �	  g	  U	  !	  	  �  �  �  |  {  =      �  �  �  �  q  S  .      �  �  �  m  @    �  �  �  �  ~  G  .    �  �  �  �  �  �  Z  (    �  �  �  k  S  2  1  0  	  �  �  �  v  \  D                                                                               map_=Map(map_1.data[::-1,::-1],map_1.meta)         map_1=Map(f[i])         g=fits.open(f[i])     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     #xcen=(xbl+xtr)*0.5;ycen=(ybl+ytr)*0.5     print 'Reading...'+f[0] def get_hmi_submap(f,xbl,ybl,xtr,ytr):       return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=Map(d[::-1,::-1],h)                 d=d[0:db.shape[0],0:db.shape[1]]-db             else:                 d=d-db[0:d.shape[0],0:d.shape[1]]             if(d.shape[0]<db.shape[0]):         else:             d=d-db         if(d.shape[0]==db.shape[0]):         h,d=aa.meta,aa.data         aa=Map(f[i])         hb,db=ab.meta,ab.data         ab=Map(f[i-1])     for i in range(1,n):     n=len(f)-1;maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] def get_hmi_rundiff_maps(f):     return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=Map(d[::-1,::-1],aa.meta)                 d=d[0:db.shape[0],0:db.shape[1]]-db             else:                 d=d-db[0:d.shape[0],0:d.shape[1]]             if(d.shape[0]<db.shape[0]):         else:             d=d-db         if(d.shape[0]==db.shape[0]):         hb,db=ab.meta,ab.data         h,d=aa.meta,aa.data         ab=Map(f[0])         aa=Map(f[i])     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] def get_hmi_basediff_maps(f): #############################################################      return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=Map(d,h)                 d=d[0:db.shape[0],0:db.shape[1]]-db             else:                 d=d-db[0:d.shape[0],0:d.shape[1]]             if(d.shape[0]<db.shape[0]):         else:             d=d-db         if(d.shape[0]==db.shape[0]):             aa=idl2sunpy_hmi(f[i]);h,d=aa.meta,aa.data             ab=idl2sunpy_hmi(f[i-1]);hb,db=ab.meta,ab.data         if(inst=='HMI'):             aa=idl2sunpy_sdo(f[i],wave,inst);h,d=aa.meta,aa.data             ab=idl2sunpy_sdo(f[i-1],wave,inst);hb,db=ab.meta,ab.data         if(inst=='AIA'):     for i in range(1,n):     n=len(f)-1;maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] def get_sunpy_rundiff_maps(f,wave,inst):       return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=Map(d,h)                 d=d[0:db.shape[0],0:db.shape[1]]-db             else:                 d=d-db[0:d.shape[0],0:d.shape[1]]             if(d.shape[0]<db.shape[0]):         else:             d=d-db         if(d.shape[0]==db.shape[0]):         hb,db=ab.meta,ab.data         h,d=aa.meta,aa.data             ab=idl2sunpy_hmi(f[0])             aa=idl2sunpy_hmi(f[i])         if(inst=='HMI'):             ab=idl2sunpy_sdo(f[0],wave,inst)             aa=idl2sunpy_sdo(f[i],wave,inst)         if(inst=='AIA'):     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] def get_sunpy_basediff_maps(f,wave,inst):      return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=Map(f[i])     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     print 'Reading...'+f[0] ad     P     G       �  E  �  �  �  �  h  P  /  .    �  �  �  s  Y     �  �  u  G  �  �  =    �
  �
  �
  �
  v
  u
  W
  D
  
  �	  ~	  }	  r	  q	  b	  P	  �  �  M  �  �  N  �  �  Q    �  �  J    �  �  9  �  �  �  x  D    �  �  p  8  �  �  P  O                              allmaps['aia171']={'map171':map171,'data171':data171,'time171':time171}     allmaps['aia131']={'map131':map131,'data131':data131,'time131':time131}     allmaps={};allmaps['aia94']={'map94':map94,'data94':data94,'time94':time94}     #map1700,data1700,time1700=get_sunpy_maps(list1700)     #map1600,data1600,time1600=get_sunpy_maps(list1600)     #map193,data193,time193=get_sunpy_maps(list193)     #map211,data211,time211=get_sunpy_maps(list211)     #map171,data171,time171=get_sunpy_maps(list171)     #map335,data335,time335=get_sunpy_maps(list335)     #map131,data131,time131=get_sunpy_maps(list131)     #map94,data94,time94=get_sunpy_maps(list94)     ################     map1700,data1700,time1700=get_sunpy_maps_rot(list1700,'1700','AIA')     map1600,data1600,time1600=get_sunpy_maps_rot(list1600,'1600','AIA')     map335,data335,time335=get_sunpy_maps_rot(list335,'335','AIA')     map304,data304,time304=get_sunpy_maps_rot(list304,'304','AIA')     map211,data211,time211=get_sunpy_maps_rot(list211,'211','AIA')     map193,data193,time193=get_sunpy_maps_rot(list193,'193','AIA')     map171,data171,time171=get_sunpy_maps_rot(list171,'171','AIA')     map131,data131,time131=get_sunpy_maps_rot(list131,'131','AIA')     map94,data94,time94=get_sunpy_maps_rot(list94,'94','AIA')     list94=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/94/*rot.sav'))     list211=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/211/*rot.sav'))     list171=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/171/*rot.sav'))     list193=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/193/*rot.sav'))     list131=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/131/*rot.sav'))     list304=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/304/*rot.sav'))     list335=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/335/*rot.sav'))     list1700=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/1700/*rot.sav'))     list1600=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/1600/*rot.sav')) if(dump_submaps): dump_submaps=1  sys.exit()      g.close()     g.writeto('/media/rohit/VLA/20160409/sun_L_20160409T1844-1846UT.50ms.cal.pol.LL.spw.0_16-31.time.18:45:10.-18:45:10.05.fits')     g[0].header['CRVAL1']=xc;g[0].header['CRVAL2']=yc     g=fits.open(f) def change_pointing(f,xc,yc):      return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=map_         maplist[i]=map_.submap(bl,tr)         tr = SkyCoord(xtr*u.arcsec, ytr*u.arcsec, frame=map_.coordinate_frame)         bl = SkyCoord(xbl*u.arcsec, ybl*u.arcsec, frame=map_.coordinate_frame)         #cent_pix=map_.world_to_pixel(SkyCoord(xcen*u.arcsec, ycen*u.arcsec, frame=map_.coordinate_frame))          map_=Map(g[0].data[0][0],g[0].header)         #g[0].data[np.isnan(g[0].data)]=0         #g[0].header['CRVAL1']=-731.12;g[0].header['CRVAL2']=243.5         #g[0].header['CRVAL1']=-770;g[0].header['CRVAL2']=220         #g[0].header['CRVAL1']=0;g[0].header['CRVAL2']=0         g=fits.open(f[i])     for i in range(n):     n=len(f);maplist=[0]*n;datalist=[0]*n;time=[0]*n     #xcen=(xbl+xtr)*0.5;ycen=(ybl+ytr)*0.5     print 'Reading...'+f[0] def get_evla_submap(f,xbl,ybl,xtr,ytr):      return maplist,datalist,time     time=np.array(time)         time[i]=produce_tstring(maplist[i])         datalist[i]=maplist[i].data         maplist[i]=map_         maplist[i]=map_.submap(bl,tr)         tr = SkyCoord(xtr*u.arcsec, ytr*u.arcsec, frame=map_.coordinate_frame)         bl = SkyCoord(xbl*u.arcsec, ybl*u.arcsec, frame=map_.coordinate_frame)         #cent_pix=map_.world_to_pixel(SkyCoord(xcen*u.arcsec, ycen*u.arcsec, frame=map_.coordinate_frame))  ad      �      7       �  h    �  }  *    �  �  �  F  �  �  h    �  �  ;  �
  �
  ?
  �	  �	  C	  �  �  @  �  �  n  O  	  �  s  (  �  �  G  �  �  N  �  �  R  �  �  V  �  �  �  )  	      �       dump_submaps=0       ###########################     pickle.dump(allmapsb,open('/media/rohit/VLA/20160409/20160409_submap_aia_base_50ms.p','wb'))     print "Writing.."     allmapsb['aiab1700']={'mapb1700':mapb1700,'datab1700':datab1700,'timeb1700':timeb1700}     allmapsb['aiab1600']={'mapb1600':mapb1600,'datab1600':datab1600,'timeb1600':timeb1600}     allmapsb['aiab335']={'mapb335':mapb335,'datab335':datab335,'timeb335':timeb335}     allmapsb['aiab304']={'mapb304':mapb304,'datab304':datab304,'timeb304':timeb304}     allmapsb['aiab211']={'mapb211':mapb211,'datab211':datab211,'timeb211':timeb211}     allmapsb['aiab193']={'mapb193':mapb193,'datab193':datab193,'timeb193':timeb193}     allmapsb['aiab171']={'mapb171':mapb171,'datab171':datab171,'timeb171':timeb171}     allmapsb['aiab131']={'mapb131':mapb131,'datab131':datab131,'timeb131':timeb131}     allmapsb={};allmapsb['aiab94']={'mapb94':mapb94,'datab94':datab94,'timeb94':timeb94}     mapb1700,datab1700,timeb1700=get_sunpy_basediff_maps(list1700,'1700','AIA')     mapb1600,datab1600,timeb1600=get_sunpy_basediff_maps(list1600,'1600','AIA')     mapb211,datab211,timeb211=get_sunpy_basediff_maps(list211,'211','AIA')     mapb193,datab193,timeb193=get_sunpy_basediff_maps(list193,'193','AIA')     mapb171,datab171,timeb171=get_sunpy_basediff_maps(list171,'171','AIA')     mapb304,datab304,timeb304=get_sunpy_basediff_maps(list304,'304','AIA')     mapb335,datab335,timeb335=get_sunpy_basediff_maps(list335,'335','AIA')     mapb131,datab131,timeb131=get_sunpy_basediff_maps(list131,'131','AIA')     mapb94,datab94,timeb94=get_sunpy_basediff_maps(list94,'94','AIA')     ##########################     pickle.dump(allmapsd,open('/media/rohit/VLA/20160409/20160409_submap_aia_diff_50ms.p','wb'))     print "Writing.."     allmapsd['aiad1700']={'mapd1700':mapd1700,'datad1700':datad1700,'timed1700':timed1700}     allmapsd['aiad1600']={'mapd1600':mapd1600,'datad1600':datad1600,'timed1600':timed1600}     allmapsd['aiad335']={'mapd335':mapd335,'datad335':datad335,'timed335':timed335}     allmapsd['aiad304']={'mapd304':mapd304,'datad304':datad304,'timed304':timed304}     allmapsd['aiad211']={'mapd211':mapd211,'datad211':datad211,'timed211':timed211}     allmapsd['aiad193']={'mapd193':mapd193,'datad193':datad193,'timed193':timed193}     allmapsd['aiad171']={'mapd171':mapd171,'datad171':datad171,'timed171':timed171}     allmapsd['aiad131']={'mapd131':mapd131,'datad131':datad131,'timed131':timed131}     allmapsd={};allmapsd['aiad94']={'mapd94':mapd94,'datad94':datad94,'timed94':timed94}     mapd1700,datad1700,timed1700=get_sunpy_rundiff_maps(list1700,'1700','AIA')     mapd1600,datad1600,timed1600=get_sunpy_rundiff_maps(list1600,'1600','AIA')     mapd193,datad193,timed193=get_sunpy_rundiff_maps(list193,'193','AIA')     mapd211,datad211,timed211=get_sunpy_rundiff_maps(list211,'211','AIA')     mapd171,datad171,timed171=get_sunpy_rundiff_maps(list171,'171','AIA')     mapd335,datad335,timed335=get_sunpy_rundiff_maps(list335,'335','AIA')     mapd304,datad304,timed304=get_sunpy_rundiff_maps(list304,'304','AIA')     mapd131,datad131,timed131=get_sunpy_rundiff_maps(list131,'131','AIA')     mapd94,datad94,timed94=get_sunpy_rundiff_maps(list94,'94','AIA')     ##########################     sys.exit()     pickle.dump(allmaps,open('/media/rohit/VLA/20160409/20160409_submap_aia_50ms.p','wb'))     print "Writing.."     allmaps['aia1700']={'map1700':map1700,'data1700':data1700,'time1700':time1700}     allmaps['aia1600']={'map1600':map1600,'data1600':data1600,'time1600':time1600}     allmaps['aia335']={'map335':map335,'data335':data335,'time335':time335}     allmaps['aia304']={'map304':map304,'data304':data304,'time304':time304}     allmaps['aia211']={'map211':map211,'data211':data211,'time211':time211}     allmaps['aia193']={'map193':map193,'data193':data193,'time193':time193} ad  &   �      ,       �  �  W  �  �  :  �  |    �  _  :  �    �
  �
  K
  �	  	  �  �  2  �  h    �  9  �  f  E  �  q  $  �  �  G    �  �  ?  �  �  y  �   �                                             allmaps={};allvlamaps0={};allvlamaps1={};allvlamaps2={};allvlamaps3={};allvlamaps4={};allvlamaps5={};allvlamaps6={};allvlamaps7={}     mapvla7,datavla7,timevla7=get_evla_submap(listvla7,0,-1,0,-1)     mapvla6,datavla6,timevla6=get_evla_submap(listvla6,0,-1,0,-1)     mapvla5,datavla5,timevla5=get_evla_submap(listvla5,0,-1,0,-1)     mapvla4,datavla4,timevla4=get_evla_submap(listvla4,0,-1,0,-1)     mapvla3,datavla3,timevla3=get_evla_submap(listvla3,0,-1,0,-1)     mapvla2,datavla2,timevla2=get_evla_submap(listvla2,0,-1,0,-1)     mapvla1,datavla1,timevla1=get_evla_submap(listvla1,0,-1,0,-1)     mapvla0,datavla0,timevla0=get_evla_submap(listvla0,0,-1,0,-1)     sys.exit()             pickle.dump(allmaps,open('/media/rohit/VLA/20160409/vlamaps_RR/vlamap_'+str(listvla0[i].split('.')[8])+'_'+"%04d"%i+'.p','wb'))             allmaps={};allmaps['vla']={'mapvla':mapvla[i],'timevla':timevla}             #allmaps={};allmaps['vla']={'mapvla':mapvla,'datavla':datavla,'timevla':timevla}             datavla[i]=datavla0[i]+datavla1[i]+datavla2[i]+datavla3[i]+datavla4[i]+datavla5[i]+datavla6[i]+datavla7[i]             print len(mapvla[i])             mapvla[i]=mapvla0[i]+mapvla1[i]+mapvla2[i]+mapvla3[i]+mapvla4[i]+mapvla5[i]+mapvla6[i]+mapvla7[i]                 mapvla7[i][k],datavla7[i][k],timevla=get_evla_submap([listvla7[i+2399*k]],0,-1,0,-1)                 mapvla6[i][k],datavla6[i][k],timevla=get_evla_submap([listvla6[i+2399*k]],0,-1,0,-1)                 mapvla5[i][k],datavla5[i][k],timevla=get_evla_submap([listvla5[i+2399*k]],0,-1,0,-1)                 mapvla4[i][k],datavla4[i][k],timevla=get_evla_submap([listvla4[i+2399*k]],0,-1,0,-1)                 mapvla3[i][k],datavla3[i][k],timevla=get_evla_submap([listvla3[i+2399*k]],0,-1,0,-1)                 mapvla2[i][k],datavla2[i][k],timevla=get_evla_submap([listvla2[i+2399*k]],0,-1,0,-1)                 mapvla1[i][k],datavla1[i][k],timevla=get_evla_submap([listvla1[i+2399*k]],0,-1,0,-1)                 mapvla0[i][k],datavla0[i][k],timevla=get_evla_submap([listvla0[i+2399*k]],0,-1,0,-1)             for k in range(4):             datavla0[i]=[0]*4;datavla1[i]=[0]*4;datavla2[i]=[0]*4;datavla3[i]=[0]*4;datavla4[i]=[0]*4;datavla5[i]=[0]*4;datavla6[i]=[0]*4;datavla7[i]=[0]*4             mapvla0[i]=[0]*4;mapvla1[i]=[0]*4;mapvla2[i]=[0]*4;mapvla3[i]=[0]*4;mapvla4[i]=[0]*4;mapvla5[i]=[0]*4;mapvla6[i]=[0]*4;mapvla7[i]=[0]*4         if(os.path.isfile('/media/rohit/VLA/20160409/vlamaps_RR/vlamap_'+str(listvla0[i].split('.')[8])+'_'+"%04d"%i+'.p')==False):         print str(listvla0[i].split('.')[8]),i     for i in range(0,2399):     datavla0=[0]*2399;datavla1=[0]*2399;datavla2=[0]*2399;datavla3=[0]*2399;datavla4=[0]*2399;datavla5=[0]*2399;datavla6=[0]*2399;datavla7=[0]*2399     mapvla0=[0]*2399;mapvla1=[0]*2399;mapvla2=[0]*2399;mapvla3=[0]*2399;mapvla4=[0]*2399;mapvla5=[0]*2399;mapvla6=[0]*2399;mapvla7=[0]*2399     mapvla=[0]*2399;datavla=[0]*2399     listvla7=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_7/*.spw.7_*FITS'))     listvla6=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_6/*.spw.6_*FITS'))     listvla5=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_5/*.spw.5_*FITS'))     listvla4=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_4/*.spw.4_*FITS'))     listvla3=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_3/*.spw.3_*FITS'))     listvla2=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_2/*.spw.2_*FITS'))     listvla1=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_1/*.spw.1_*FITS'))     listvla0=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_0/*.spw.0_*FITS'))     #listvla=sorted(glob.glob('/media/rohit/VLA/20160409/images_1s/sun*FITS'))     #mapvla,datavla,timevla=get_evla_submap(listvla,-1000,100,-600,400) if(dump_submaps): ad     ,     C       �  Q     �  Q  �  �  D  �  �  D  �  �  7  �
  �
  �
  r
  H
  4
  &
  %
  
  
  
  
  �	  �	  �	  �	  �	  m	  l	  [	  G	  �  �  i  Q  �  �  �  �  �  j  ?    �  �  Z  "  �  �  �  �  Q    �  �  @  �  �  #  �  '  �  ,                      maxTbv[i][j]=[0]*2000;xcvmax[i][j]=[0]*2000;ycvmax[i][j]=[0]*2000;Tbv_r1[i][j]=[0]*2000;Tbv_r2[i][j]=[0]*2000             listvla_v=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_V/spw_'+str(i)+'/*spw.*'+spc[j]+'*.FITS'))[0:2000]             maxTbi[i][j]=[0]*2000;xcimax[i][j]=[0]*2000;ycimax[i][j]=[0]*2000;Tbi_r1[i][j]=[0]*2000;Tbi_r2[i][j]=[0]*2000             listvla_r=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_'+str(i)+'/*spw.*'+spc[j]+'*.FITS'))[0:2000]             listvla_l=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_LL/spw_'+str(i)+'/*spw.*'+spc[j]+'*.FITS'))[0:2000]         for j in range(4):         xci90[i]=[0]*4;yci90[i]=[0]*4;xcv90[i]=[0]*4;ycv90[i]=[0]*4;xcl90[i]=[0]*4;ycl90[i]=[0]*4;xcr90[i]=[0]*4;ycr90[i]=[0]*4         Tbl_r1[i]=[0]*4;Tbl_r2[i]=[0]*4;Tbr_r1[i]=[0]*4;Tbr_r2[i]=[0]*4;areai50[i]=[0]*4         Tbi_r1[i]=[0]*4;Tbi_r2[i]=[0]*4;Tbv_r1[i]=[0]*4;Tbv_r2[i]=[0]*4         maxTbr[i]=[0]*4;xcrmax[i]=[0]*4;ycrmax[i]=[0]*4         maxTbl[i]=[0]*4;xclmax[i]=[0]*4;yclmax[i]=[0]*4         maxTbi[i]=[0]*4;xcimax[i]=[0]*4;ycimax[i]=[0]*4         maxTbv[i]=[0]*4;xcvmax[i]=[0]*4;ycvmax[i]=[0]*4     for i in range(8):     areai50=[0]*8     Tbl_r1=[0]*8;Tbl_r2=[0]*8;Tbr_r1=[0]*8;Tbr_r2=[0]*8     Tbi_r1=[0]*8;Tbi_r2=[0]*8;Tbv_r1=[0]*8;Tbv_r2=[0]*8     xci90=[0]*8;yci90=[0]*8;xcv90=[0]*8;ycv90=[0]*8;xcl90=[0]*8;ycl90=[0]*8;xcr90=[0]*8;ycr90=[0]*8     maxTbr=[0]*8;xcrmax=[0]*8;ycrmax=[0]*8     maxTbl=[0]*8;xclmax=[0]*8;yclmax=[0]*8     maxTbi=[0]*8;xcimax=[0]*8;ycimax=[0]*8     maxTbv=[0]*8;xcvmax=[0]*8;ycvmax=[0]*8     spc=['0-15','16-31','32-47','48-63'] if(get_max): get_max=1          mapvla_i[k],datavla_i[k],timevla=get_evla_submap([listvla_i[k]],0,-1,0,-1)         mapvla_v[k],datavla_v[k],timevla=get_evla_submap([listvla_v[k]],0,-1,0,-1)     for k in range(32):     mapvla_v=[0]*32;datavla_v=[0]*32;mapvla_i=[0]*32;datavla_i=[0]*32     listvla_i=sorted(glob.glob('/media/rohit/VLA/20160409/images_I/*FITS'))     listvla_v=sorted(glob.glob('/media/rohit/VLA/20160409/images_V/*FITS')) if(get_submap_pol): get_submap_pol=1  ################ Only radio analysis   gtime=goes['tarray'] gflux=goes['yclean'] goes=readsav('/media/rohit/VLA/20160409/20160409_idlsave_goes.sav')  ################ GOES  sys.exit()      return mi     mi=Map(nd,meta)     meta=ml.meta;nd=(ml.data+mr.data)*0.5 def get_mapI(ml,mr):      pickle.dump(allvlamaps7,open('/media/rohit/VLA/20160409/20160409_vla_spw_7_50ms.p','wb'))     allvlamaps7['vla7']={'mapvla':mapvla7,'datavla':datavla7,'timevla':timevla7}     pickle.dump(allvlamaps6,open('/media/rohit/VLA/20160409/20160409_vla_spw_6_50ms.p','wb'))     allvlamaps6['vla6']={'mapvla':mapvla6,'datavla':datavla6,'timevla':timevla6}     pickle.dump(allvlamaps5,open('/media/rohit/VLA/20160409/20160409_vla_spw_5_50ms.p','wb'))     allvlamaps5['vla5']={'mapvla':mapvla5,'datavla':datavla5,'timevla':timevla5}     pickle.dump(allvlamaps4,open('/media/rohit/VLA/20160409/20160409_vla_spw_4_50ms.p','wb'))     allvlamaps4['vla4']={'mapvla':mapvla4,'datavla':datavla4,'timevla':timevla4}     pickle.dump(allvlamaps3,open('/media/rohit/VLA/20160409/20160409_vla_spw_3_50ms.p','wb'))     allvlamaps3['vla3']={'mapvla':mapvla3,'datavla':datavla3,'timevla':timevla3}     pickle.dump(allvlamaps2,open('/media/rohit/VLA/20160409/20160409_vla_spw_2_50ms.p','wb'))     allvlamaps2['vla2']={'mapvla':mapvla2,'datavla':datavla2,'timevla':timevla2}     pickle.dump(allvlamaps1,open('/media/rohit/VLA/20160409/20160409_vla_spw_1_50ms.p','wb'))     allvlamaps1['vla1']={'mapvla':mapvla1,'datavla':datavla1,'timevla':timevla1}     pickle.dump(allvlamaps0,open('/media/rohit/VLA/20160409/20160409_vla_spw_0_50ms.p','wb'))     allvlamaps0['vla0']={'mapvla':mapvla0,'datavla':datavla0,'timevla':timevla0} ad  1        1       �  �  A    �  �  w  .  �  �    �  P    �
  �
  C
  �	  �	  o	  W	  	  �  r  �  �  \  /     �    �  �  �  t  �  �    �  �  �    �  �  m  3  �  �                                                                       ycrmax[i][j][k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xcrmax[i][j][k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 yc,xc=np.where(Tbr==np.nanmax(Tbr))                 Tbr=h.data;maxTbr[i][j][k]=np.nanmax(Tbr)                 h=mr[0]                 #######                 ycl90[i][j][k]=h.reference_coordinate.Ty.value+(ycf-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xcl90[i][j][k]=h.reference_coordinate.Tx.value+(xcf-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 xcf,ycf=ut.fitEllipse(bi)[0:2]                 bi=ut.get_bimage(Tbl_f,0.95)                 Tbl_f=Tbl*1.0;Tbl_f[np.isnan(Tbl_f)]=0                 Tbl_r1[i][j][k]=Tbl[138:148,120:130].mean();Tbl_r2[i][j][k]=Tbl[124:136,116:126].mean()                 yclmax[i][j][k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xclmax[i][j][k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 yc,xc=np.where(Tbl==np.nanmax(Tbl))                 Tbl=h.data;maxTbl[i][j][k]=np.nanmax(Tbl)                 h=ml[0]                 #######                 ycv90[i][j][k]=h.reference_coordinate.Ty.value+(ycf-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xcv90[i][j][k]=h.reference_coordinate.Tx.value+(xcf-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 xcf,ycf=ut.fitEllipse(bi)[0:2]                 bi=ut.get_bimage(Tbv_f,0.95)                 Tbv_f=Tbv*1.0;Tbv_f[np.isnan(Tbv_f)]=0                 Tbv_r1[i][j][k]=Tbv[138:148,120:130].mean();Tbv_r2[i][j][k]=Tbv[124:136,116:126].mean()                 ycvmax[i][j][k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xcvmax[i][j][k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 yc,xc=np.where(Tbv==np.nanmax(Tbv))                 Tbv=h.data;maxTbv[i][j][k]=np.nanmax(Tbv)                 h=mv[0]                 mv,dv,tv=get_evla_submap([listvla_v[k]],0,-1,0,-1)                 ######                 yci90[i][j][k]=hl.reference_coordinate.Ty.value+(ycf-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value                 xci90[i][j][k]=hl.reference_coordinate.Tx.value+(xcf-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value                 xcf,ycf=ut.fitEllipse(bi)[0:2]                 bi=ut.get_bimage(Tbi_f,0.95)                 Tbi_f=Tbi*1.0;Tbi_f[np.isnan(Tbi_f)]=0                 areai50[i][j][k]=len(np.where(Tbi>np.nanmax(Tbi)*0.5)[0])*2.0                 Tbi_r1[i][j][k]=Tbi[138:148,120:130].mean();Tbi_r2[i][j][k]=Tbi[124:136,116:126].mean()                 ycimax[i][j][k]=hl.reference_coordinate.Ty.value+(yc-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value                 xcimax[i][j][k]=hl.reference_coordinate.Tx.value+(xc-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value                 yc,xc=np.where(Tbi==np.nanmax(Tbi))                 Tbi=(hl.data+hr.data)*0.5;maxTbi[i][j][k]=np.nanmax(Tbi)                 hl=ml[0];hr=mr[0]                 mr,dr,tr=get_evla_submap([listvla_r[k]],0,-1,0,-1)                 ml,dl,tl=get_evla_submap([listvla_l[k]],0,-1,0,-1)             for k in range(2000):             xci90[i][j]=[0]*2000;yci90[i][j]=[0]*2000;xcv90[i][j]=[0]*2000;ycv90[i][j]=[0]*2000;xcl90[i][j]=[0]*2000;ycl90[i][j]=[0]*2000;xcr90[i][j]=[0]*2000;ycr90[i][j]=[0]*2000             maxTbr[i][j]=[0]*2000;xcrmax[i][j]=[0]*2000;ycrmax[i][j]=[0]*2000;Tbr_r1[i][j]=[0]*2000;Tbr_r2[i][j]=[0]*2000;areai50[i][j]=[0]*2000             maxTbl[i][j]=[0]*2000;xclmax[i][j]=[0]*2000;yclmax[i][j]=[0]*2000;Tbl_r1[i][j]=[0]*2000;Tbl_r2[i][j]=[0]*2000 ad  -        4       �  a  4    �    �  �  +  �  W  �  �  H    �
  R
  
  �	  �	  f	  �  �  x  =    �  O    �  �  c  (  �  �  �  <    �  W  �  s  N      �  �  x    �  3                                                       for k in range(2000):     mapvla_v=[0]*2000;datavla_v=[0]*2000;mapvla_i=[0]*2000;datavla_i=[0]*2000;timevla=[0]*2000;mapvla_l=[0]*2000;mapvla_r=[0]*2000     listvla_rr=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_RR/spw_0/*FITS'))[0:2000]     listvla_ll=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_LL/spw_0/*FITS'))[0:2000]     listvla_v=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_V/spw_0/*spw.0_16*.FITS'))[0:2000] if(get_submap_pol): get_submap_pol=1  #Tbmayn[np.where(ycmax<255)]=np.nan;Tbmays[np.where(ycmax>255)]=np.nan #Tbmayn=maxTbi*1.0;Tbmays=maxTbi*1.0 xcrmax,ycrmax,xcr90,ycr90,maxTbr,Tbr_r1,Tbr_r2=pickle.load(open('/media/rohit/VLA/20160409/vlamax_loc_r.p','rb')) xclmax,yclmax,xcl90,ycl90,maxTbl,Tbl_r1,Tbl_r2=pickle.load(open('/media/rohit/VLA/20160409/vlamax_loc_l.p','rb')) xcimax,ycimax,xci90,yci90,maxTbi,Tbi_r1,Tbi_r2,areai50=pickle.load(open('/media/rohit/VLA/20160409/vlamax_loc_i.p','rb')) #Tbmayn[np.where(ycmax<255)]=np.nan;Tbmays[np.where(ycmax>255)]=np.nan Tbmayn=maxTbv*1.0;Tbmays=maxTbv*1.0 xcvmax,ycvmax,xcv90,ycv90,maxTbv,Tbv_r1,Tbv_r2=pickle.load(open('/media/rohit/VLA/20160409/vlamax_loc_v.p','rb'))       pickle.dump([xcrmax,ycrmax,xcr90,ycr90,maxTbr,Tbr_r1,Tbr_r2],open('/media/rohit/VLA/20160409/vlamax_loc_r.p','wb'))     Tbr_r2=np.array(Tbr_r2);Tbr_r2=Tbr_r2.reshape(32,2000)     Tbr_r1=np.array(Tbr_r1);Tbr_r1=Tbr_r1.reshape(32,2000)     ycrmax=np.array(ycrmax);ycrmax=ycrmax.reshape(32,2000)     xcrmax=np.array(xcrmax);xcrmax=xcrmax.reshape(32,2000)     maxTbr=np.array(maxTbr);maxTbr=maxTbr.reshape(32,2000)     pickle.dump([xclmax,yclmax,xcl90,ycl90,maxTbl,Tbl_r1,Tbl_r2],open('/media/rohit/VLA/20160409/vlamax_loc_l.p','wb'))     Tbl_r2=np.array(Tbl_r2);Tbl_r2=Tbl_r2.reshape(32,2000)     Tbl_r1=np.array(Tbl_r1);Tbl_r1=Tbl_r1.reshape(32,2000)     yclmax=np.array(yclmax);yclmax=yclmax.reshape(32,2000)     xclmax=np.array(xclmax);xclmax=xclmax.reshape(32,2000)     maxTbl=np.array(maxTbl);maxTbl=maxTbl.reshape(32,2000)     pickle.dump([xcvmax,ycvmax,xcv90,ycv90,maxTbv,Tbv_r1,Tbv_r2],open('/media/rohit/VLA/20160409/vlamax_loc_v.p','wb'))     Tbv_r2=np.array(Tbv_r2);Tbv_r2=Tbv_r2.reshape(32,2000)     Tbv_r1=np.array(Tbv_r1);Tbv_r1=Tbv_r1.reshape(32,2000)     ycvmax=np.array(ycvmax);ycvmax=ycvmax.reshape(32,2000)     xcvmax=np.array(xcvmax);xcvmax=xcvmax.reshape(32,2000)     maxTbv=np.array(maxTbv);maxTbv=maxTbv.reshape(32,2000)     pickle.dump([xcimax,ycimax,xci90,yci90,maxTbi,Tbi_r1,Tbi_r2,areai50],open('/media/rohit/VLA/20160409/vlamax_loc_i.p','wb'))     Tbi_r2=np.array(Tbi_r2);Tbi_r2=Tbi_r2.reshape(32,2000)     Tbi_r1=np.array(Tbi_r1);Tbi_r1=Tbi_r1.reshape(32,2000)     xcr90=np.array(xcr90);xcr90=xcr90.reshape(32,2000);ycr90=np.array(ycr90);ycr90=ycr90.reshape(32,2000)     xcl90=np.array(xcl90);xcl90=xcl90.reshape(32,2000);ycl90=np.array(ycl90);ycl90=ycl90.reshape(32,2000)     xcv90=np.array(xcv90);xcv90=xcv90.reshape(32,2000);ycv90=np.array(ycv90);ycv90=ycv90.reshape(32,2000)     xci90=np.array(xci90);xci90=xci90.reshape(32,2000);yci90=np.array(yci90);yci90=yci90.reshape(32,2000)     xcimax=np.array(xcimax);xcimax=xcimax.reshape(32,2000);ycimax=np.array(ycimax);ycimax=ycimax.reshape(32,2000)     maxTbi=np.array(maxTbi);maxTbi=maxTbi.reshape(32,2000)     areai50=np.array(areai50);areai50=areai50.reshape(32,2000)                 ycr90[i][j][k]=h.reference_coordinate.Ty.value+(ycf-(h.reference_pixel.y.value-1))*h.scale.axis2.value                 xcr90[i][j][k]=h.reference_coordinate.Tx.value+(xcf-(h.reference_pixel.x.value-1))*h.scale.axis1.value                 xcf,ycf=ut.fitEllipse(bi)[0:2]                 bi=ut.get_bimage(Tbr_f,0.95)                 Tbr_f=Tbr*1.0;Tbr_f[np.isnan(Tbr_f)]=0                 Tbr_r1[i][j][k]=Tbr[138:148,120:130].mean();Tbr_r2[i][j][k]=Tbr[124:136,116:126].mean() ad     Z     I       �  p  6    �  �  �  �  �  C  �  f  E    �  �  �  0  �  p  0    �
  �
  G
  �	  H	  �  2  �  �  �  �  [  <  �  �  v  6  5  �  �  �  �  p  o  _  B    �  �  �  6  �  �  �  `  _  )    �  �  T    �  �  �  �  �  �  �  w  Z  Y                                ax1.plot(gtime,gflux[1])     ax1.plot(gtime,gflux[0])     f,(ax1,ax2,ax3)=plt.subplots(3,1,figsize=(15,15)) if(plot_ds): plot_ds=1    b_proj_euv = utils.skycoord_to_pixel(b_hp_euv, pmap.wcs) b_proj_ls = utils.skycoord_to_pixel(b_hp_ls, pmap.wcs) b_proj_fr = utils.skycoord_to_pixel(b_hp_fr, pmap.wcs) from astropy.wcs import utils b_hp_fr,b_hp_ls,b_hp_euv,hmiwcs=pickle.load(open('/media/rohit/VLA/paraview/bproj.p','rb')) pmap=allmaps['aia171']['map171'][0] ######################## Extrapolated Magnetic Fields  freq=np.round(np.linspace(0.994,2.006,32),3) dx_km=1400 mapex_by=pickle.load(open('/media/rohit/VLA/20160409_EUV/20160409_by.p','rb')) mapex_bx=pickle.load(open('/media/rohit/VLA/20160409_EUV/20160409_bx.p','rb')) mapex_bz=pickle.load(open('/media/rohit/VLA/20160409_EUV/20160409_bz.p','rb')) mapex_babs=pickle.load(open('/media/rohit/VLA/20160409_EUV/20160409_babs.p','rb')) from astropy.wcs import WCS from astropy.coordinates import SkyCoord from sunpy.coordinates import frames from scipy.io import readsav # Extrapolation  hmimap=Map(hmid,hmimap.meta) hmid[np.where(hmid<-5000)]=0 hmid=hmimap.data[::-1,::-1] hmimap=Map(hmifile) hmifile='/media/rohit/VLA/20160409_EUV/hmi.m_45s.2016.04.09_18_45_00_TAI.magnetogram.fits'  maphmir,datalistr,time=get_sunpy_rundiff_maps(hmilist,'','HMI') maphmib,datalistb,time=get_sunpy_basediff_maps(hmilist,'','HMI') maphmi,datahmi,timehmi=get_sunpy_maps_rot(hmilist,'','HMI') #    maphmi[k],datahmi[k],timevla=get_hmi_submap([hmilist[k]],0,-1,0,-1) #for k in range(len(hmilist)): maphmi=[0]*len(hmilist);datahmi=[0]*len(hmilist) hmilist=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/hmi/*rot.sav')) ############### HMI  timevla_all1=np.hstack((np.array(qstimevla)[:,0],timevla_all))  TbLLr1,TbLLr2,TbLLr3,TbLLr4,TbLLr5,xcLLmax,ycLLmax,xcLL90,ycLL90,timevla_all=pickle.load(open('/media/rohit/VLA/20160409/MaxLL.p','rb')) qsx,qsy,qsxcr90,qsycr90,qsmaxTbr,qsTbr_r1,qsTbr_r2,qsarear50,qstimevla=pickle.load(open('/media/rohit/VLA/20160409/vlamax_loc_r_qs.p','rb'))     pickle.dump([xcrmax,ycrmax,qsxcr90,qsycr90,maxTbr,Tbr_r1,Tbr_r2,arear50,qstimevla],open('/media/rohit/VLA/20160409/vlamax_loc_r_qs.p','wb'))         qsycr90[k]=hl.reference_coordinate.Ty.value+(ycf-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value         qsxcr90[k]=hl.reference_coordinate.Tx.value+(xcf-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value         xcf,ycf=ut.fitEllipse(bi)[0:2]         bi=ut.get_bimage(Tbr_f,0.95)         Tbr_f=Tbr*1.0;Tbr_f[np.isnan(Tbr_f)]=0         arear50[k]=len(np.where(Tbr>np.nanmax(Tbr)*0.5)[0])*2.0         Tbr_r1[k]=Tbr[138:148,120:130].mean();Tbr_r2[k]=Tbr[124:136,116:126].mean()         ycrmax[k]=hl.reference_coordinate.Ty.value+(yc-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value         xcrmax[k]=hl.reference_coordinate.Tx.value+(xc-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value         yc,xc=np.where(Tbr==np.nanmax(Tbr))         Tbr=hl.data;maxTbr[k]=np.nanmax(Tbr)         hl=m[0]         m,d,qstimevla[k]=get_evla_submap([listqs[k]],0,-1,0,-1)     for k in range(len(listqs)):     qsxcr90=[0]*len(listqs);qsycr90=[0]*len(listqs)     xcrmax=[0]*len(listqs);ycrmax=[0]*len(listqs);maxTbr=[0]*len(listqs);Tbr_r1=[0]*len(listqs);Tbr_r2=[0]*len(listqs);arear50=[0]*len(listqs);qstimevla=[0]*len(listqs)     listqs=sorted(glob.glob('/media/rohit/VLA/20160409/1844/fits_0_16-31/*spw.0*FITS')) if(get_qs): get_qs=1  vlamax_v=np.nanmax(np.array(datavla_v),axis=(1,2,3))         mapvla_l[k]=ml;mapvla_r[k]=mr         mapvla_i[k]=get_mapI(ml[0],mr[0])         mr,d,t=get_evla_submap([listvla_rr[k]],0,-1,0,-1)         ml,d,t=get_evla_submap([listvla_ll[k]],0,-1,0,-1)         mapvla_v[k],datavla_v[k],timevla[k]=get_evla_submap([listvla_v[k]],0,-1,0,-1) ad  t   x     :       �  �  �  �  �  �  �  �  i    �  c    �  �  �  �  �  r  L  +  N    �  �  A    �
  �
  �	  �	  �  \  �  E  �  �  m    �  {  g  f  X  G  /  	  �    �  i  Q  �  �  �  F  �  x  w                                                                                                                              dd0=Map(dcp_data,mapvla_i[i][0].meta)         dcp_data=mapvla_v[i][0].data*100/mapvla_i[i][0].data;dcp_data[np.isnan(dcp_data)]=0;dcp_data[np.where(dcp_data<0)]=0;dcp_data[np.where(dcp_data>100)]=0         lev2=np.array([1,5,10,20,50,60,70,80,90])*u.percent         lev1=np.array([10,20,30,40,50,60,70,80,90])*u.percent         lev0=np.array([50,55,60,65,70,75,80,85,90])*u.percent         #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent         #cc.draw_grid()         p=hmimap.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-2000,vmax=2000)         xlaia=-1037.6;xraia=1031.6;ylaia=-1031.2;yraia=1031.9         #xlaia=cc.center.Tx.value-0.6*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.6*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.6*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.6*int(cc.data.shape[0]/2)         ax0 = f.add_subplot(111)         f=plt.figure(figsize=(10,10))     for i in range(32): if(plot_vi_hmi): plot_vi_hmi=1          plt.close()         plt.savefig('pngs_dcp_hmi/dcp_hmi_'+"%02d"%i+'.png')         ax0.text(-840,330,'Contours (%): 50, 55, 60, 65, 70, 75, 80, 85, 90',color='yellow')         ax0.text(-840,210,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='blue')         ax0.set_xlim([-850,-700]);ax0.set_ylim([200,350])         #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])         #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')         #mapvla_v[i][0].draw_contours(levels=lev1,colors='yellow',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         #mapvla_i[i][0].draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)         dd0=Map(dcp_data,mapvla_i[i][0].meta)         dcp_data=mapvla_v[i][0].data*100/mapvla_i[i][0].data;dcp_data[np.isnan(dcp_data)]=0;dcp_data[np.where(dcp_data<0)]=0;dcp_data[np.where(dcp_data>100)]=0         lev2=np.array([1,5,10,20,50,60,70,80,90])*u.percent         lev1=np.array([10,20,30,40,50,60,70,80,90])*u.percent         lev0=np.array([50,55,60,65,70,75,80,85,90])*u.percent         #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent         #cc.draw_grid()         p=hmimap.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-2000,vmax=2000)         xlaia=-1037.6;xraia=1031.6;ylaia=-1031.2;yraia=1031.9         #xlaia=cc.center.Tx.value-0.6*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.6*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.6*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.6*int(cc.data.shape[0]/2)         ax0 = f.add_subplot(111)         f=plt.figure(figsize=(10,10))     for i in range(32): if(plot_dcp_hmi): plot_dcp_hmi=1      plt.close()     plt.savefig('/media/rohit/VLA/20160409/spec_max/max_poss_'+"%02d"%i+'.png')     ax.legend();ax.set_title(str(freq[i])+' GHz');ax.set_ylim(0,40);ax.set_xlim(0,100)     ax.set_ylabel('$T_B$ (MK)');ax.set_ylabel('$T_B$ (MK)');ax.set_xlabel('Time (sec)')     ax.plot(np.arange(2000)*0.05,Tbmays[i]/1.e6,'o',color='red',label='South Source')     #ax.plot(np.arange(2000)*0.05,Tbmayn[i]/1.e6,'o',color='blue',label='North Source')     f,ax=plt.subplots(1,1,figsize=(15,6)) for i in range(32): i=0 plot_position=1        plt.show()     ax2.imshow(TbLLr1.swapaxes(0,1),aspect='auto') ad          7         �  .  �    �  {  A  �  �  Y  E  D  6  %    �
  �
  L
  =
  <
  ;
  0
  "
  

  �	  �	  ]	  ,	  O    �  �  d  &  �  �    �  �  ~    �  �  �  Y    �  j  )                             plot_dcp=1            plt.close()         plt.savefig('pngs_vi_aia171/vi_aia171_'+"%02d"%i+'.png')         ax0.text(-840,330,'Contours (%): 50, 55, 60, 65, 70, 75, 80, 85, 90',color='yellow')         ax0.text(-840,210,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='blue')         ax0.set_xlim([-850,-700]);ax0.set_ylim([200,350])         #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])         #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')         mapvla_v[i][0].draw_contours(levels=lev1,colors='yellow',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i][0].draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i][0].data[np.isnan(mapvla_i[i][0].data)]=0;mapvla_v[i][0].data[np.isnan(mapvla_v[i][0].data)]=0         #dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)         dd0=Map(dcp_data,mapvla_i[i][0].meta)         dcp_data=mapvla_v[i][0].data*100/mapvla_i[i][0].data;dcp_data[np.isnan(dcp_data)]=0;dcp_data[np.where(dcp_data<0)]=0;dcp_data[np.where(dcp_data>100)]=0         lev2=np.array([1,5,10,20,50,60,70,80,90])*u.percent         lev1=np.array([10,20,30,40,50,60,70,80,90])*u.percent         lev0=np.array([50,55,60,65,70,75,80,85,90])*u.percent         #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent         #cc.draw_grid()         p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=-1230;xraia=-569;ylaia=-47.9;yraia=572         #xlaia=cc.center.Tx.value-0.6*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.6*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.6*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.6*int(cc.data.shape[0]/2)         cc=allmaps['aia171']['map171'][tidx_171]         tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],allmaps['aia171']['time171'][0])[0]         ax0 = f.add_subplot(111)         f=plt.figure(figsize=(10,10))     for i in range(32): if(plot_dcp): plot_dcp=1       plt.show()     ax0.set_ylabel('DCP (%)');ax0.set_xlabel('Frequency (GHz)')     ax0.plot(freq,maxTbv[:,770:870].mean(axis=1)/maxTbi[:,770:870].mean(axis=1)*100,'o-')     ax0 = f.add_subplot(111)     f=plt.figure(figsize=(10,10)) if(plot_dcp_2d): plot_dcp_2d=1          plt.close()         plt.savefig('pngs_vi_hmi/vi_hmi_'+"%02d"%i+'.png')         ax0.text(-840,330,'Contours (%): 10,20,30,40,50,60,70,80,90',color='yellow')         ax0.text(-840,210,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='blue')         ax0.set_xlim([-850,-700]);ax0.set_ylim([200,350])         #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])         #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')         mapvla_v[i][0].draw_contours(levels=lev1,colors='yellow',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i][0].draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i][0].data[np.isnan(mapvla_i[i][0].data)]=0;mapvla_v[i][0].data[np.isnan(mapvla_v[i][0].data)]=0         #dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2) ad     �      1       �  �  �  E    7    �  �  L    �  �  �  �  �
  >
  �	  J	  �  a     �  �  1  �  B  .  -  ,  !    �  �  �  G    �  �  �  �  p  %  �  �  ]  �  �  �   �                            dcp_data=mapvla_v[i][0].data*100/mapvla_i[i].data*(mapvla_v[i][0].data/np.nanmax(mapvla_v[i][0].data));dcp_data[np.isnan(dcp_data)]=0;dcp_data[np.where(dcp_data<0)]=0;dcp_data[np.where(dcp_data>100)]=0         lev2=np.array([1,5,10,20,50,60,70,80,90])*u.percent         lev1=np.array([30,40,50,60,70,80,90])/np.nanmax(mapvla_v[i][0].data)*(4.e7)*u.percent         #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent         #cc.draw_grid()         #p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-80,vmax=80)         p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=-1230;xraia=-569;ylaia=-47.9;yraia=572         #xlaia=cc.center.Tx.value-0.6*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.6*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.6*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.6*int(cc.data.shape[0]/2)         #cc=Map(cc0.data-cc1.data,cc0.meta)         #cc1=allmaps['aia171']['map171'][tidx_171-1]         #cc0=allmaps['aia171']['map171'][tidx_171]         cc=allmaps['aia171']['map171'][tidx_171]         tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],timevla[i])[0]         f,ax=plt.subplots(2,1,figsize=(8,15));ax0=ax[0];ax1=ax[1]     for i in range(800,1200):     #for i in range(2000): if(plot_dcp): plot_dcp=1           plt.close()         plt.savefig('pngs_v_aia171_time/dcp_aia171_'+"%02d"%i+'.png')         ax1.plot(np.arange(2000)*0.05,vlamax_v,'-',label='Stokes V');ax1.axvline(x=i*0.05,color='k');ax1.set_xlabel('Time (sec)');ax1.set_ylabel('T$_{B}$');ax1.legend()         ax0.text(-840,330,'Contours (%): 50, 55, 60, 65, 70, 75, 80, 85, 90',color='yellow')         ax0.text(-840,210,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='blue')         ax0.set_xlim([-850,-700]);ax0.set_ylim([200,350])         #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])         #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')         #mapvla_v[i][0].draw_contours(levels=lev1,colors='yellow',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         #mapvla_i[i].draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i].data[np.isnan(mapvla_i[i].data)]=0;mapvla_v[i][0].data[np.isnan(mapvla_v[i][0].data)]=0         dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)         dd0=Map(dcp_data,mapvla_i[i].meta)         dcp_data=mapvla_v[i][0].data*100/mapvla_i[i].data*(mapvla_v[i][0].data/np.nanmax(mapvla_v[i][0].data));dcp_data[np.isnan(dcp_data)]=0;dcp_data[np.where(dcp_data<0)]=0;dcp_data[np.where(dcp_data>100)]=0         lev2=np.array([1,5,10,20,50,60,70,80,90])*u.percent         lev1=np.array([30,40,50,60,70,80,90])*u.percent         lev0=np.array([50,55,60,65,70,75,80,85,90])*u.percent         #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent         #cc.draw_grid()         p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')         xlaia=-1230;xraia=-569;ylaia=-47.9;yraia=572         #xlaia=cc.center.Tx.value-0.6*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.6*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.6*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.6*int(cc.data.shape[0]/2)         cc=allmaps['aia171']['map171'][tidx_171]         tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],timevla[i])[0]         f,ax=plt.subplots(2,1,figsize=(8,15));ax0=ax[0];ax1=ax[1]     for i in range(2000): if(plot_dcp): ad  F   Z     >       �    �    �  +  �  C    �  p    �
  
  �	  �	  \	  H	  G	  F	  &	  	  �  �  �  �  f  F  &    �  �  �  �  ?  �  �  X  �  �  �  �  �  9  �  �  �  �    �  ^  2  �  �  �  �  x    �  �  �  Z  Y                                                                            yc,xc=np.where(Tbl==np.nanmax(Tbl))     Tbl=hl.data     hl=mapvla_l[k][0]     ycimed[k]=hi.reference_coordinate.Ty.value+(yc-(hi.reference_pixel.y.value-1))*hi.scale.axis2.value     xcimed[k]=hi.reference_coordinate.Tx.value+(xc-(hi.reference_pixel.x.value-1))*hi.scale.axis1.value         yc,xc=idx[0][1],idx[0][0]     else:         yc,xc=idx[1],idx[0]     if(len(idx[0])==1):     idx=np.where(np.abs(Tbi-np.nanmedian(Tbi))==np.nanmin(np.abs(Tbi-np.nanmedian(Tbi))))     Tbi[np.where(Tbi<Tbi.max()*0.5)]=np.nan     Tbi_r1[k]=hi.data[124:137,121:124].mean();Tbi_r2[k]=hi.data[138:141,123:126].mean()     ycimax[k]=hi.reference_coordinate.Ty.value+(yc-(hi.reference_pixel.y.value-1))*hi.scale.axis2.value     xcimax[k]=hi.reference_coordinate.Tx.value+(xc-(hi.reference_pixel.x.value-1))*hi.scale.axis1.value     yc,xc=np.where(Tbi==np.nanmax(Tbi))     Tbi=hi.data     hi=mapvla_i[k][0]     ycvmed[k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value     xcvmed[k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value         yc,xc=idx[0][1],idx[0][0]     else:         yc,xc=idx[1],idx[0]     if(len(idx[0])==1):     idx=np.where(np.abs(Tbv-np.nanmedian(Tbv))==np.nanmin(np.abs(Tbv-np.nanmedian(Tbv))))     Tbv[np.where(Tbv<Tbv.max()*0.5)]=np.nan     Tbv_r1[k]=h.data[124:137,121:124].mean();Tbv_r2[k]=h.data[138:141,123:126].mean()     ycvmax[k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value     xcvmax[k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value     yc,xc=np.where(Tbv==np.nanmax(Tbv))     Tbv=h.data     h=mapvla_v[k][0] for k in range(2000): Tbr_r1=[0]*2000;Tbr_r2=[0]*2000 Tbl_r1=[0]*2000;Tbl_r2=[0]*2000 Tbv_r1=[0]*2000;Tbv_r2=[0]*2000 Tbi_r1=[0]*2000;Tbi_r2=[0]*2000 xcimed=[0]*2000;ycimed=[0]*2000 xcimax=[0]*2000;ycimax=[0]*2000 xcvmed=[0]*2000;ycvmed=[0]*2000 xcrmax=[0]*2000;ycrmax=[0]*2000 xclmax=[0]*2000;yclmax=[0]*2000 xcvmax=[0]*2000;ycvmax=[0]*2000           plt.close()         plt.savefig('pngs_v_aia171_time/v_abs_aia171_'+"%02d"%i+'.png')         #plt.savefig('pngs_v_aia171_time/dcp_run_aia171_'+"%02d"%i+'.png')         ax1.set_xlim(40,60)         ax1.plot(np.arange(2000)*0.05,vlamax_v,'o-',label='Stokes V');ax1.axvline(x=i*0.05,color='k');ax1.set_xlabel('Time (sec)');ax1.set_ylabel('T$_{B}$');ax1.legend()         ax0.text(-840,330,'Contours (%): 20, 22, 24, 26, 28, 30, 32, 34, 36 MK',color='green')         #ax0.text(-840,330,'Contours (%): 50, 55, 60, 65, 70, 75, 80, 85, 90',color='blue')         ax0.text(-840,210,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='blue')         ax0.set_xlim([-850,-700]);ax0.set_ylim([200,350])         #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])         #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')         mapvla_v[i][0].draw_contours(levels=lev1,colors='yellow',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         #mapvla_i[i].draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         mapvla_i[i].data[np.isnan(mapvla_i[i].data)]=0;mapvla_v[i][0].data[np.isnan(mapvla_v[i][0].data)]=0         #dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])         xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)         lev0=np.array([50,55,60,65,70,75,80,85,90])/100*np.nanmax(dd0.data)*u.percent         dd0=Map(dcp_data,mapvla_i[i].meta) ad  -   A     >       �  0  �  �  �  �  "  �  b  ]  \  [  W  C  �  �  D  �  x    �
  �
  �
  �
  �
  V
  
  �	  ,	  �  \  �  �  �  �  �  z  <  �  �  R  �  ~  #  �  I  9  8  �  �  ]  �  �  �  �  N  "  �  �  M  B  A  @                                                plt.show() ax1.set_ylabel('$T_B$ (MK)');ax0.set_ylabel('Y-Coordinate (arcsec)');ax1.set_xlabel('Time (sec)') ax1.plot(np.arange(len(y))*0.05,np.hstack((qsTbr_r1,Tbr_r1[1]))/1.e6,'o-') ax0.plot(np.arange(len(y))*0.05,y,'o-') y=np.hstack((np.array(qsy)[:,0],ycrmax[1])) f,ax=plt.subplots(2,1,figsize=(8,15),sharex=True);ax0=ax[0];ax1=ax[1]  plt.show() ax1.set_ylabel('$T_B$ (MK)');ax0.set_ylabel('T$_B$ (MK)');ax1.set_xlabel('Time (sec)') ax1.plot(np.arange(2000)*0.05,(np.array(Tb_r2)-np.array(Tb_r1))/1.e6,'o-',label='R2-R1');ax1.legend() ax0.plot(np.arange(2000)*0.05,np.array(Tb_r2)/1.e6,'o-',label='R2');ax0.legend() ax0.plot(np.arange(2000)*0.05,np.array(Tb_r1)/1.e6,'o-',label='R1') f,ax=plt.subplots(2,1,figsize=(8,15),sharex=True);ax0=ax[0];ax1=ax[1]      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_spec/dcp_spec_regions_'+"%02d"%i+'.png')     ax1.set_ylabel('DCP (V/I) (\%)');ax0.set_ylabel('T$_b$ (MK)');ax0.set_xlabel('time (sec)');ax1.set_xlabel('Frequency (MHz)')     ax1.set_ylim(0,100);ax0.set_ylim(0,50);ax0.legend();ax0.set_title(str(freq[0])+' GHz')     ax1.plot(freq,(np.array(Tbv_r2[:,i])/np.array(Tbi_r2[:,i]))*100,'o-',label='R2 (South)');ax1.legend()     ax1.plot(freq,(np.array(Tbv_r1[:,i])/np.array(Tbi_r1[:,i]))*100,'o-',label='R1 (North)');ax1.legend()     ax0.axvline(x=np.arange(2000)[i]*0.05,color='k')     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r2[0])/1.e6,'-',label='R2 (South)');ax0.legend()     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r1[0])/1.e6,'-',label='R1 (North)') #     f,ax=plt.subplots(2,1,figsize=(15,8));ax0=ax[0];ax1=ax[1] for i in range(2000): i=0      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_spec/Tbi_dcp_regions_'+"%02d"%i+'.png')     ax1.set_ylabel('DCP (V/I) (\%)');ax0.set_ylabel('T$_b$ (MK)');ax1.set_xlabel('time (sec)')     ax1.set_ylim(0,100);ax0.set_ylim(0,50);ax0.legend();ax0.set_title(str(freq[i])+' GHz')     ax1.plot(np.arange(2000)*0.05,(np.array(Tbv_r2[i])/np.array(Tbi_r2[i]))*100,'-',label='R2 (South)');ax1.legend()     ax1.plot(np.arange(2000)*0.05,(np.array(Tbv_r1[i])/np.array(Tbi_r1[i]))*100,'-',label='R1 (North)');ax1.legend()     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r2[i])/1.e6,'-',label='R2 (South)');ax0.legend()     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r1[i])/1.e6,'-',label='R1 (North)') #     f,ax=plt.subplots(2,1,figsize=(15,8),sharex=True);ax0=ax[0];ax1=ax[1] for i in range(32): i=0      plt.close()     plt.savefig('/media/rohit/VLA/20160409/pngs_spec/Tbi_regions_'+"%02d"%i+'.png')     ax1.set_ylabel('$T_B$ (MK)');ax0.set_ylabel('T$_B$ (MK)');ax1.set_xlabel('time (sec)')     ax1.set_ylim(-8,12);ax0.set_ylim(0,50);ax0.legend();ax0.set_title(str(freq[i])+' GHz')     ax1.plot(np.arange(2000)*0.05,(np.array(Tbi_r2[i])-np.array(Tbi_r1[i]))/1.e6,'-',label='R2-R1');ax1.legend()     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r2[i])/1.e6,'-',label='R2 (South)');ax0.legend()     ax0.plot(np.arange(2000)*0.05,np.array(Tbi_r1[i])/1.e6,'-',label='R1 (North)') #     f,ax=plt.subplots(2,1,figsize=(15,8),sharex=True);ax0=ax[0];ax1=ax[1] for i in range(32): i=0            Tbr_r1[k]=hi.data[124:137,121:124].mean();Tbr_r2[k]=hi.data[138:141,123:126].mean()     yclmax[k]=hl.reference_coordinate.Ty.value+(yc-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value     xclmax[k]=hl.reference_coordinate.Tx.value+(xc-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value     yc,xc=np.where(Tbl==np.nanmax(Tbl))     Tbr=hr.data     hr=mapvla_r[k][0]     Tbl_r1[k]=hl.data[124:137,121:124].mean();Tbl_r2[k]=hl.data[138:141,123:126].mean()     yclmax[k]=hl.reference_coordinate.Ty.value+(yc-(hl.reference_pixel.y.value-1))*hl.scale.axis2.value     xclmax[k]=hl.reference_coordinate.Tx.value+(xc-(hl.reference_pixel.x.value-1))*hl.scale.axis1.value ad  #   W     F       �  �  ]  �  �  �  �  q  Z  �  �  \  4  �  d  Y  X  A    �  �    �
  �
  �
  a
  1
  
  �	  �	  d	  +	  �  Z  -     �  �  y  J    �  �  �  �  �  x  =    �  I  -  �  �  �  m  =    �  �  g  *  �  i  <    �  �  �  W  V                                     ax1.plot(t[1153],vlamax_v[1153],'o',color='r') ax1.plot(t[1058],vlamax_v[1058],'o',color='g') ax1.plot(t[966],vlamax_v[966],'o',color='r') ax1.plot(t[954],vlamax_v[954],'o',color='r') ax1.plot(t[883],vlamax_v[883],'o',color='g') ax1.plot(t[858],vlamax_v[858],'o',color='g') ax1.plot(t[781],vlamax_v[781],'o',color='g') ax1.plot(t,vlamax_v,'o-',label='Stokes V');ax1.axvline(x=i*0.05,color='k');ax1.set_xlabel('Time (sec)');ax1.set_ylabel('T$_{B}$');ax1.legend(loc=4) #ax0.plot(xcvmax[1057:1062],ycvmax[1057:1062],'o',color='g') #ax0.plot(xcvmax[944:950],ycvmax[944:950],'o',color='r') #ax0.plot(xcvmax[880:885],ycvmax[880:885],'o',color='g') ax0.plot(xcvmax[1153],ycvmax[1153],'o',color='r') ax0.plot(xcvmax[1058],ycvmax[1058],'o',color='g') ax0.plot(xcvmax[966],ycvmax[966],'o',color='r') ax0.plot(xcvmax[954],ycvmax[954],'o',color='r') ax0.plot(xcvmax[883],ycvmax[883],'o',color='g') ax0.plot(xcvmax[858],ycvmax[858],'o',color='g') ax0.plot(xcvmax[781],ycvmax[781],'o',color='g') f.colorbar(p,label='B (G)') xlaia=-949;xraia=-649.1;ylaia=70;yraia=369.4;p=mapex_bz[0].plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-750,vmax=750) #p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') #cc=allmaps['aia171']['map171'][20] f,ax=plt.subplots(2,1,figsize=(12,15));ax0=ax[0];ax1=ax[1] t=np.arange(2000)*0.05  plt.show() ax1.set_xlim(35,60) #ax1.plot(t[964:970],vlamax_v[964:970],'o',color='r') #ax1.plot(t[855:860],vlamax_v[855:860],'o',color='g') ax1.plot(t[1153],vlamax_v[1153],'o',color='r') ax1.plot(t[1058],vlamax_v[1058],'o',color='g') ax1.plot(t[966],vlamax_v[966],'o',color='r') ax1.plot(t[954],vlamax_v[954],'o',color='r') ax1.plot(t[883],vlamax_v[883],'o',color='g') ax1.plot(t[858],vlamax_v[858],'o',color='g') ax1.plot(t[781],vlamax_v[781],'o',color='g') ax1.plot(t,vlamax_v,'o-',label='Stokes V');ax1.axvline(x=i*0.05,color='k');ax1.set_xlabel('Time (sec)');ax1.set_ylabel('T$_{B}$');ax1.legend(loc=4) #ax0.plot(xcvmax[1057:1062],ycvmax[1057:1062],'o',color='g') #ax0.plot(xcvmax[944:950],ycvmax[944:950],'o',color='r') #ax0.plot(xcvmax[880:885],ycvmax[880:885],'o',color='g') ax0.plot(xcvmax[1153],ycvmax[1153],'o',color='r') ax0.plot(xcvmax[1058],ycvmax[1058],'o',color='g') ax0.plot(xcvmax[966],ycvmax[966],'o',color='r') ax0.plot(xcvmax[954],ycvmax[954],'o',color='r') ax0.plot(xcvmax[883],ycvmax[883],'o',color='g') ax0.plot(xcvmax[858],ycvmax[858],'o',color='g') ax0.plot(xcvmax[781],ycvmax[781],'o',color='g') f.colorbar(p,label='B (G)') xlaia=-1037.6;xraia=1031.6;ylaia=-1031.2;yraia=1031.9;p=hmimap.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',vmin=-2000,vmax=2000) #p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') #cc=allmaps['aia171']['map171'][20] f,ax=plt.subplots(2,1,figsize=(8,15));ax0=ax[0];ax1=ax[1] t=np.arange(2000)*0.05  plt.show() ax1.set_ylabel('$T_B$ (MK)');ax0.set_ylabel('Y-Coordinate (arcsec)');ax1.set_xlabel('Time (sec)') ax1.plot(t1,vlamax_v1/1.e6,'o',markersize=8,color='r');ax1.plot(t2,vlamax_v2/1.e6,'o',markersize=8,color='g') ax1.plot(t,vlamax_v/1.e6,'-',color='k') ax0.plot(t1,ycvmax1,'o',color='r');ax0.plot(t2,ycvmax2,'o',color='g') f,ax=plt.subplots(2,1,figsize=(8,15),sharex=True);ax0=ax[0];ax1=ax[1] t1=t[idx1];ycvmax1=ycvmax[idx1];t2=t[idx2];ycvmax2=ycvmax[idx2];vlamax_v1=vlamax_v[idx1];vlamax_v2=vlamax_v[idx2] t=np.arange(2000)*0.05 idx1=np.where(ycvmax<255)[0];idx2=np.where(ycvmax>255)[0] ycvmax=np.array(ycvmax).flatten();xcvmax=np.array(xcvmax).flatten()  plt.show() ax1.set_ylabel('$T_B$ (MK)');ax0.set_ylabel('Y-Coordinate (arcsec)');ax1.set_xlabel('Time (sec)') ax1.plot(np.arange(2000)*0.05,vlamax_v/1.e6,'o-') ax0.plot(np.arange(2000)*0.05,ycvmax,'o-') f,ax=plt.subplots(2,1,figsize=(8,15),sharex=True);ax0=ax[0];ax1=ax[1] ad  J   Z     =       �  �  �  u  t  )  �  �    �      �  {    �
  �
  g
  c
  K
  '
  �	  ^	  N	  6	  	  �  �  �  �  q    �  g  �  �  B  �  �  a        
    �  �  +      �  �  �  �  e  >  �  d  4  �  Z  Y                                                                                    ycRRmax[v][k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value         xcRRmax[v][k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value         yc,xc=np.where(TbRRv==np.nanmax(TbRRv))         ycRR90[v][k]=h.reference_coordinate.Ty.value+(ycf-(h.reference_pixel.y.value-1))*h.scale.axis2.value         xcRR90[v][k]=h.reference_coordinate.Tx.value+(xcf-(h.reference_pixel.x.value-1))*h.scale.axis1.value         xcf,ycf=ut.fitEllipse(bi)[0:2]         bi=ut.get_bimage(TbRRv_f,0.95)         TbRRv_f[np.isnan(TbRRv_f)]=0         TbRRv_f=TbRRv*1.0         TbRRv=h.data         h=d['vla']['mapvla'][k][0]     for k in range(32):     print vfile     TbRRr1[v]=[0]*32;TbRRr2[v]=[0]*32;TbRRr3[v]=[0]*32;TbRRr4[v]=[0]*32;TbRRr5[v]=[0]*32;xcRRmax[v]=[0]*32;ycRRmax[v]=[0]*32;xcRR90[v]=[0]*32;ycRR90[v]=[0]*32     d=pickle.load(open(vfile,'rb')) for vfile in vlalistRR: v=0       v=v+1         TbLLr5[v][k]=np.nanmax(TbLLv[re[4][0]:re[4][1],re[4][2]:re[4][3]])         TbLLr4[v][k]=np.nanmax(TbLLv[re[3][0]:re[3][1],re[3][2]:re[3][3]])         TbLLr3[v][k]=np.nanmax(TbLLv[re[2][0]:re[2][1],re[2][2]:re[2][3]])         TbLLr2[v][k]=np.nanmax(TbLLv[re[1][0]:re[1][1],re[1][2]:re[1][3]])         TbLLr1[v][k]=np.nanmax(TbLLv[re[0][0]:re[0][1],re[0][2]:re[0][3]])         ycLLmax[v][k]=h.reference_coordinate.Ty.value+(yc-(h.reference_pixel.y.value-1))*h.scale.axis2.value         xcLLmax[v][k]=h.reference_coordinate.Tx.value+(xc-(h.reference_pixel.x.value-1))*h.scale.axis1.value         yc,xc=np.where(TbLLv==np.nanmax(TbLLv))         ycLL90[v][k]=h.reference_coordinate.Ty.value+(ycf-(h.reference_pixel.y.value-1))*h.scale.axis2.value         xcLL90[v][k]=h.reference_coordinate.Tx.value+(xcf-(h.reference_pixel.x.value-1))*h.scale.axis1.value         xcf,ycf=ut.fitEllipse(bi)[0:2]         bi=ut.get_bimage(TbLLv_f,0.95)         TbLLv_f[np.isnan(TbLLv_f)]=0         TbLLv_f=TbLLv*1.0         TbLLv=h.data         h=d['vla']['mapvla'][k][0]     for k in range(32):     print vfile     TbLLr1[v]=[0]*32;TbLLr2[v]=[0]*32;TbLLr3[v]=[0]*32;TbLLr4[v]=[0]*32;TbLLr5[v]=[0]*32;xcLLmax[v]=[0]*32;ycLLmax[v]=[0]*32;xcLL90[v]=[0]*32;ycLL90[v]=[0]*32     timevla_all[v]=d['vla']['timevla'][0]     d=pickle.load(open(vfile,'rb')) for vfile in vlalistLL: v=0 freq=np.linspace(0.994,2.006,32) timevla_all=[0]*len(vlalistLL) xcRR90=[0]*len(vlalistRR);ycRR90=[0]*len(vlalistRR);xcLL90=[0]*len(vlalistLL);ycLL90=[0]*len(vlalistLL) xcRRmax=[0]*len(vlalistRR);ycRRmax=[0]*len(vlalistRR);xcLLmax=[0]*len(vlalistLL);ycLLmax=[0]*len(vlalistLL) ycRRr1=[0]*len(vlalistRR);ycRRr2=[0]*len(vlalistRR);ycRRr3=[0]*len(vlalistRR);ycRRr4=[0]*len(vlalistRR);ycRRr5=[0]*len(vlalistRR) xcRRr1=[0]*len(vlalistRR);xcRRr2=[0]*len(vlalistRR);xcRRr3=[0]*len(vlalistRR);xcRRr4=[0]*len(vlalistRR);xcRRr5=[0]*len(vlalistRR) TbRRr1=[0]*len(vlalistRR);TbRRr2=[0]*len(vlalistRR);TbRRr3=[0]*len(vlalistRR);TbRRr4=[0]*len(vlalistRR);TbRRr5=[0]*len(vlalistRR) ycLLr1=[0]*len(vlalistLL);ycLLr2=[0]*len(vlalistLL);ycLLr3=[0]*len(vlalistLL);ycLLr4=[0]*len(vlalistLL);ycLLr5=[0]*len(vlalistLL) xcLLr1=[0]*len(vlalistLL);xcLLr2=[0]*len(vlalistLL);xcLLr3=[0]*len(vlalistLL);xcLLr4=[0]*len(vlalistLL);xcLLr5=[0]*len(vlalistLL) TbLLr1=[0]*len(vlalistLL);TbLLr2=[0]*len(vlalistLL);TbLLr3=[0]*len(vlalistLL);TbLLr4=[0]*len(vlalistLL);TbLLr5=[0]*len(vlalistLL) re=[[124,134,120,130],[140,150,90,100],[95,115,70,90],[105,125,30,50],[95,115,95,115]] vlalistRR=sorted(glob.glob('/media/rohit/VLA/20160409/vlamaps_RR/vla*.p')) vlalistLL=sorted(glob.glob('/media/rohit/VLA/20160409/vlamaps_LL/vla*.p'))  plt.show() ax1.set_xlim(35,60) #ax1.plot(t[964:970],vlamax_v[964:970],'o',color='r') #ax1.plot(t[855:860],vlamax_v[855:860],'o',color='g') ad     E     C       �  j    �  �      �  �  �  �  U  �  �  �  �  g  �
  �
  �
  �
  {
  l
  
  �	  b	  D	  9	  8	  	  �  �  +  �  �  �  �  �  t  �  �  E    �  �  �  �  h  >    �  �  w  g  \  [  Z  "    �  _    �  %  �  s  E  D                               ax[0,1].text(25,25,' Region 5',color='white') ax[0,0].text(25,25,' Region 1',color='white') ax[0,0].set_xlabel('Time (sec)');ax[1,0].set_xlabel('Time (sec)');ax[0,1].set_xlabel('Time (sec)');ax[1,1].set_xlabel('Time (sec)') ax[0,0].set_ylabel('Frequency (GHz)');ax[1,0].set_ylabel('Frequency (GHz)');ax[0,1].set_ylabel('Frequency (GHz)');ax[1,1].set_ylabel('Frequency (GHz)') ax[1,1].imshow(TbLLr4.swapaxes(0,1),aspect='auto',origin=0,vmin=1.e6,vmax=10.e6) ax[0,1].imshow(TbLLr3.swapaxes(0,1),aspect='auto',origin=0,vmin=1.e6,vmax=10.e6) ax[1,0].imshow(TbLLr5.swapaxes(0,1),aspect='auto',origin=0,vmin=1.e6,vmax=10.e6) im1=ax[0,0].imshow(TbLLr1.swapaxes(0,1),aspect='auto',origin=0,vmin=1.e6,vmax=10.e6) fig, ax = plt.subplots(2, 2) from mpl_toolkits.axes_grid1 import make_axes_locatable   plt.show()     plt.close()     plt.savefig('pngs_dcp/dcp_'+"%02d"%ff+'_zoom.png')     plt.title('Frequency: '+str(np.round(freq[ff],3))+' GHz')     ax[2].set_ylim(0,50);ax[2].set_xlim(40,80)     ax[2].set_xlabel('Time (sec)')     ax[2].set_ylabel('Position (arcsec)')     ax[2].plot(x,loc_diff_LR,'o-')     ax[1].set_ylim(0,1.0)     ax[1].set_ylabel('Stokes (V/I)')     ax[1].plot(x,dcp_r1[:,ff],'o-')     ax[0].legend();ax[0].set_ylim(0,150)     ax[0].set_ylabel('Stokes I $\ T_B$ (MK)')     ax[0].plot(x,(TbLLr1[:,ff]+TbRRr1[:,ff])/1.e6,'o-',label=str(np.round(freq[ff],3))+' GHz')     fig,ax=plt.subplots(3,1,sharex=True,figsize=(10,13))     loc_diff_LR=np.sqrt((np.concatenate(xcLLmax[:,ff])[:2399]-xcRRmax[:2399,ff,0])**2 + (np.concatenate(ycLLmax[:,ff])[:2399]-ycRRmax[:2399,ff,0])**2) for ff in range(32): x=np.linspace(0,120,2399)  plt.show() ax.legend();ax1.legend(loc=2) ax.set_xlabel('Time (sec)');ax.set_ylabel('X-Centroid (arcsec)');ax1.set_ylabel('T$_B$ (MK)') ax.plot(np.linspace(0,120,2399),xcRR90.mean(axis=1)-xcLL90.mean(axis=1),'o-',color='red',label='X-Centroid (RR-LL)') ax1.plot(np.linspace(0,120,2399),TbRRr1[:,0]/1.e6,'o-',color='black',label='T$_B$') ax1=ax.twinx() fig,ax=plt.subplots(1,1,sharex=True,figsize=(10,10))  plt.show() ax.legend();ax1.legend(loc=2) ax.set_xlabel('Time (sec)');ax.set_ylabel('Y-Centroid (arcsec)');ax1.set_ylabel('T$_B$ (MK)') ax.plot(np.linspace(0,120,2399),ycRR90.std(axis=1),'o-',color='red',label='Y-Centroid') ax1.plot(np.linspace(0,120,2399),TbRRr1[:,0]/1.e6,'o-',color='black',label='T$_B$') ax1=ax.twinx() fig,ax=plt.subplots(1,1,sharex=True,figsize=(10,10))  ff=11 dcp_r1=(TbRRr1-TbLLr1)/(TbLLr1+TbRRr1) TbLLr1,TbLLr2,TbLLr3,TbLLr4,TbLLr5,xcLLmax,ycLLmax,xcLL90,ycLL90,timevla_all=pickle.load(open('/media/rohit/VLA/20160409/MaxLL.p','rb')) TbRRr1,TbRRr2,TbRRr3,TbRRr4,TbRRr5,xcRRmax,ycRRmax,xcRR90,ycRR90=pickle.load(open('/media/rohit/VLA/20160409/MaxRR.p','rb'))  #### READ  pickle.dump([TbRRr1,TbRRr2,TbRRr3,TbRRr4,TbRRr5,xcRRmax,ycRRmax,xcRR90,ycRR90],open('MaxRR.p','wb')) pickle.dump([TbLLr1,TbLLr2,TbLLr3,TbLLr4,TbLLr5,xcLLmax,ycLLmax,xcLL90,ycLL90,timevla_all],open('MaxLL.p','wb'))  xcRR90=np.array(xcRR90);ycRR90=np.array(ycRR90) xcRRmax=np.array(xcRRmax);ycRRmax=np.array(ycRRmax);xcLLmax=np.array(xcLLmax);ycLLmax=np.array(ycLLmax);xcLL90=np.array(xcLL90);ycLL90=np.array(ycLL90) TbRRr1=np.array(TbRRr1);TbRRr2=np.array(TbRRr2);TbRRr3=np.array(TbRRr3);TbRRr4=np.array(TbRRr4);TbRRr5=np.array(TbRRr5) TbLLr1=np.array(TbLLr1);TbLLr2=np.array(TbLLr2);TbLLr3=np.array(TbLLr3);TbLLr4=np.array(TbLLr4);TbLLr5=np.array(TbLLr5)     v=v+1         TbRRr5[v][k]=np.nanmax(TbRRv[re[4][0]:re[4][1],re[4][2]:re[4][3]])         TbRRr4[v][k]=np.nanmax(TbRRv[re[3][0]:re[3][1],re[3][2]:re[3][3]])         TbRRr3[v][k]=np.nanmax(TbRRv[re[2][0]:re[2][1],re[2][2]:re[2][3]])         TbRRr2[v][k]=np.nanmax(TbRRv[re[1][0]:re[1][1],re[1][2]:re[1][3]])         TbRRr1[v][k]=np.nanmax(TbRRv[re[0][0]:re[0][1],re[0][2]:re[0][3]]) ad  V   R     8       �  �  <  �  l    �  *  �  P  )  �  �  �  �  �  |  {  p  ]  H  .  �
  �
  �
  �
  �
  �
  f
  9
  
  �	  �	  �	  Y	  }  6  �  �  �  �  6    �  �  �  ,  �  �  d  �  �  9  �  o  R  Q                                                                                            ax1 = f.add_subplot(212)     ax0.add_patch(patches.Rectangle((-831,175),40,40,linewidth=5,edgecolor='magenta',facecolor='none'))     ax0.add_patch(patches.Rectangle((-961,195),40,40,linewidth=5,edgecolor='b',facecolor='none'))     ax0.add_patch(patches.Rectangle((-881,175),40,40,linewidth=5,edgecolor='red',facecolor='none'))     ax0.add_patch(patches.Rectangle((-841,265),20,20,linewidth=5,edgecolor='g',facecolor='none'))     ax0.add_patch(patches.Rectangle((-781,233),40,40,linewidth=5,edgecolor='cyan',facecolor='none'))     ax0.text(-1000,60,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='white')     ax0.set_xlim([-1000,-700]);ax0.set_ylim([50,400])     #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd1.draw_contours(levels=lev1,colors='b',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd1.center.Tx.value-2.0*int(dd1.data.shape[0]/2);xrvla=dd1.center.Tx.value+2.0*int(dd1.data.shape[0]/2);ylvla=dd1.center.Ty.value-2.0*int(dd1.data.shape[1]/2);yrvla=dd1.center.Ty.value+2.0*int(dd1.data.shape[0]/2)     dd1=vmRR;dd1.data[np.isnan(dd1.data)]=0     lev1=np.array([40,50,60,70,90])*u.percent     dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)     dd0=vmLL;dd0.data[np.isnan(dd0.data)]=0     lev0=np.array([40,50,60,70,90])*u.percent     #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     cc=allmaps['aia171']['map171'][tidx_171]     tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],timevla_all[i])[0]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(6,10))     vmRR=dRR['vla']['mapvla'][0][0]     dRR=pickle.load(open(vlalistRR[i],'rb'))     vmLL=dLL['vla']['mapvla'][0][0]     dLL=pickle.load(open(vlalistLL[i],'rb')) for i in range(2399):   Tb_r=np.array(Tb_r)         Tb_r[i][j]=np.mean(Tb1[0][j][re[i][0]:re[i][1],re[i][2]:re[i][3]])     for j in range(2399):     Tb_r[i]=[0]*2399 for i in range(5): Tb_r=[0]*5  plt.plot(TbRRr1[860],'o-') plt.plot(TbLLr1[860],'o-')  plt.show() fig.colorbar(im1, cax=cax, orientation='vertical') cax = divider.append_axes('right', size='5%', pad=0.05) divider = make_axes_locatable(ax[0,0]) ax[1,1].set_yticks(np.arange(32)[::4]);ax[1,1].set_yticklabels(np.round(np.linspace(0.994,2.006,32)[::4],2)) ax[0,1].set_yticks(np.arange(32)[::4]);ax[0,1].set_yticklabels(np.round(np.linspace(0.994,2.006,32)[::4],2)) ax[1,0].set_yticks(np.arange(32)[::4]);ax[1,0].set_yticklabels(np.round(np.linspace(0.994,2.006,32)[::4],2)) ax[0,0].set_yticks(np.arange(32)[::4]);ax[0,0].set_yticklabels(np.round(np.linspace(0.994,2.006,32)[::4],2)) ax[1,1].set_xticks([0,480,960,1440,1920,2400]);ax[1,1].set_xticklabels(['0','24','48','72','98','120']) ax[1,0].set_xticks([0,480,960,1440,1920,2400]);ax[1,0].set_xticklabels(['0','24','48','72','98','120']) ax[0,1].set_xticks([0,480,960,1440,1920,2400]);ax[0,1].set_xticklabels(['0','24','48','72','98','120']) ax[0,0].set_xticks([0,480,960,1440,1920,2400]);ax[0,0].set_xticklabels(['0','24','48','72','98','120']) ax[1,1].text(25,25,' Region 4',color='white') ax[1,0].text(25,25,' Region 3',color='white') ad  .        4       �  Q  �  �  J  �  �  B  �  �  ^  !  �  �  �  �  �  z  g  ]  0    �
  �
  �
  }
  ,
  �	  #	  �  �  _  3  S  �  �  �  �  &  �  �  Z    �  <  �  t    �  �  Y                                                        ax1.set_yscale('linear');ax1.set_ylim(0,50);ax1.grid(True)     ax1.legend(fontsize=10)#;ax1.set_ylim(0,100)     ax1.plot(Tbi_r1[0:8].mean(axis=0)/1.e6,'o-',markersize=2,label='Region 1 (Stokes-I)',color='k')     ax1 = f.add_subplot(212)     #ax0.add_patch(patches.Rectangle((-831,175),40,40,linewidth=5,edgecolor='magenta',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-961,195),40,40,linewidth=5,edgecolor='b',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-881,175),40,40,linewidth=5,edgecolor='red',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-841,265),20,20,linewidth=5,edgecolor='g',facecolor='none'))     #ax0.add_patch(patches.Rectangle((-781,233),40,40,linewidth=5,edgecolor='cyan',facecolor='none'))     ax0.text(-1000,60,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='white')     ax0.set_xlim([-900,-700]);ax0.set_ylim([150,350])     #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd1.draw_contours(levels=lev1,colors='white',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd1.center.Tx.value-2.0*int(dd1.data.shape[0]/2);xrvla=dd1.center.Tx.value+2.0*int(dd1.data.shape[0]/2);ylvla=dd1.center.Ty.value-2.0*int(dd1.data.shape[1]/2);yrvla=dd1.center.Ty.value+2.0*int(dd1.data.shape[0]/2)     dd1=vmRR;dd1.data[np.isnan(dd1.data)]=0     lev1=np.array([40,50,60,70,90])*u.percent     #dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)     dd0=vmLL;dd0.data[np.isnan(dd0.data)]=0     lev0=np.array([40,50,60,70,90])*u.percent     #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     cc=allmaps['aia171']['map171'][tidx_171]     tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],timevla_all[i])[0]     ax0 = f.add_subplot(211)     f=plt.figure(figsize=(6,10))     vmRR=dRR['vla']['mapvla'][0][0]     dRR=pickle.load(open(vlalistRR[i],'rb'))     vmLL=dLL['vla']['mapvla'][0][0]     dLL=pickle.load(open(vlalistLL[i],'rb'))     i=860 for i in range(1): #for i in range(2399):       plt.close()     plt.savefig('pngs_spec_movie/aia171_'+"%02d"%i+'.png')     ax1.set_xlabel('Frequency (GHz)');ax1.set_ylabel('$T_B$ (MK)')     ax1.set_yscale('log');ax1.set_ylim(0,300);ax1.grid(True)     ax1.legend(fontsize=10)#;ax1.set_ylim(0,100)     ax1.plot(freq,TbRRr5[i]/1.e6,'o--',markersize=2,label='Region 5 (RR)',color='magenta')     ax1.plot(freq,TbRRr4[i]/1.e6,'o--',markersize=2,label='Region 4 (RR)',color='blue')     ax1.plot(freq,TbRRr3[i]/1.e6,'o--',markersize=2,label='Region 3 (RR)',color='red')     ax1.plot(freq,TbRRr2[i]/1.e6,'o--',markersize=2,label='Region 2 (RR)',color='green')     ax1.plot(freq,TbRRr1[i]/1.e6,'o--',markersize=2,label='Region 1 (RR)',color='cyan')     ax1.plot(freq,TbLLr5[i]/1.e6,'o-',markersize=2,label='Region 5 (LL)',color='magenta')     ax1.plot(freq,TbLLr4[i]/1.e6,'o-',markersize=2,label='Region 4 (LL)',color='blue')     ax1.plot(freq,TbLLr3[i]/1.e6,'o-',markersize=2,label='Region 3 (LL)',color='red')     ax1.plot(freq,TbLLr2[i]/1.e6,'o-',markersize=2,label='Region 2 (LL)',color='green')     ax1.plot(freq,TbLLr1[i]/1.e6,'o-',markersize=2,label='Region 1 (LL)',color='cyan') ad           ;       �  Q      �  �  |  ,  �  �  �  �  �  �  �  p  (  �  �  :  �  �  /  �
  �
  �
  �
  �
  �
  S
  w	  0	  �  �  o  �    �  �  �  O  �  �  f  1  !  �  s  r  E  �  �  E  �  �  �  c  &        for i in range(len(list171)):     timstr_1600[i]= list1600[i].split('T')[-1].split('Z')[0] for i in range(len(list1600)):     timstr_vla[i]=listvla[i].split('time.')[1].split('.FITS')[0].split('-')[0] for i in range(len(listvla)): timstr_vla=[0]*len(listvla);timstr_1600=[0]*len(list1600);timstr_171=[0]*len(list171) list171=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/171/*fits')) list1600=sorted(glob.glob('/media/rohit/VLA/20160409_EUV/full_sun/1600/*fits')) listvla=sorted(glob.glob('/media/rohit/VLA/20160409/images_50ms_LL/spw_0/sun*.spw.0_16-31*FITS')) ################ Make Time String ##########      #ax0.text(-1200,50,'Contours: 20%, 30%, 40%, 50%, 60%, 70%, 80%, 90%',color='yellow')     #ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow')     plt.close()     plt.savefig('pngs_spec/aia171_'+"%02d"%i+'.png')     ax0.text(-1200,0,str(np.round(dd0.meta['crval3']/1.e9,4))+' GHz',color='green')     ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia])     #ax0.set_title('AIA 171 $\AA$:'+timstr_171[tidx171[i]]+' VLA: '+timstr_vla[i]+' UT')     dd1.draw_contours(levels=lev1,colors='b',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd1.center.Tx.value-2.0*int(dd1.data.shape[0]/2);xrvla=dd1.center.Tx.value+2.0*int(dd1.data.shape[0]/2);ylvla=dd1.center.Ty.value-2.0*int(dd1.data.shape[1]/2);yrvla=dd1.center.Ty.value+2.0*int(dd1.data.shape[0]/2)     dd1=vlaRR['vla']['mapvla'][i][0];dd1.data[np.isnan(dd1.data)]=0     lev1=np.array([40,50,60,70,90])*u.percent     dd0.draw_contours(levels=lev0,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix])     xlvla=dd0.center.Tx.value-2.0*int(dd0.data.shape[0]/2);xrvla=dd0.center.Tx.value+2.0*int(dd0.data.shape[0]/2);ylvla=dd0.center.Ty.value-2.0*int(dd0.data.shape[1]/2);yrvla=dd0.center.Ty.value+2.0*int(dd0.data.shape[0]/2)     dd0=vlaLL['vla']['mapvla'][i][0];dd0.data[np.isnan(dd0.data)]=0     lev0=np.array([40,50,60,70,90])*u.percent     #lev1=(1.5e7/dd0.data.max())*np.array([20,30,40,50,60,70,80,90])*u.percent     p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto')     xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2)     cc=allmaps['aia171']['map171'][tidx_171]     ax0 = f.add_subplot(111)     f=plt.figure(figsize=(6,6)) for i in range(32):   tidx_1600=ut.find_predecessor(allmaps['aia1600']['time1600'],vlaLL['vla']['timevla'][0])[0] tidx_193=ut.find_predecessor(allmaps['aia193']['time193'],vlaLL['vla']['timevla'][0])[0] tidx_171=ut.find_predecessor(allmaps['aia171']['time171'],vlaLL['vla']['timevla'][0])[0] tidx_131=ut.find_predecessor(allmaps['aia131']['time131'],vlaLL['vla']['timevla'][0])[0] tidx_94=ut.find_predecessor(allmaps['aia94']['time94'],vlaLL['vla']['timevla'][0])[0] vlaLL=pickle.load(open(vlafileLL,'rb'));vlaRR=pickle.load(open(vlafileRR,'rb')) vlafileRR='/media/rohit/VLA/20160409/vlamaps_RR/vlamap_18:44:43_0860.p' vlafileLL='/media/rohit/VLA/20160409/vlamaps_LL/vlamap_18:44:43_0860.p' #################  sys.exit()       plt.show()     plt.xlabel('Time (HH:MM:SS UT)');plt.ylabel('Frequency (GHz)')     plt.yticks([0,4,8,12,15],[freq[0],freq[4],freq[8],freq[12],freq[15]])     plt.xticks([0,600,1200,1800],['18:44:00','18:44:30','18:45:00','18:45:30'])     plt.colorbar(label='$T_B$ (MK)')     plt.imshow(Tbi_r1[0:16]/1.e6,aspect='auto',origin=0,cmap='YlOrRd')     plt.figure(figsize=(5,5))     plt.show()     #plt.savefig('pngs_spec_movie/aia171_'+"%02d"%i+'.png')     ax1.set_xlabel('Time (HH:MM:SS UT)');ax1.set_ylabel('$T_B$ (MK)')     ax1.set_xticks([0,600,1200,1800]);ax1.set_xticklabels(['18:44:00','18:44:30','18:45:00','18:45:30']) ad     0     ?       �  �  �  �  �  :  �  �  ?  �  �  }  (  �  �    _  �  ~  
  �
  l
  ?
  �	  �	  �	  C	  	  �  �  G  	  �  �  �  p  G      �  c    �  d    �  P  �  �  -  �  �  s        �  �  �  �  y  W  0  /                                  vlasize[k][i]=[0]*Tb0.shape[1]     for i in range(Tb0.shape[0]):     vlasize_fwhm[k]=[0]*Tb0.shape[0]     vlasize[k]=[0]*Tb0.shape[0] for k in range(len(lev)): vlasize_fwhm=[0]*len(lev) vlasize=[0]*len(lev) lev=[0.5,0.6,0.7,0.9]  vlafreqidx=np.array(list(np.arange(1))*2399).reshape(2399,1).swapaxes(0,1).flatten() #vlafreqidx=np.array(list(np.arange(32))*119).reshape(119,32).swapaxes(0,1).flatten()      #tidx1700[i]=ut.find_predecessor(allmaps['aia1700']['time1700'],vla0['vla0']['timevla'][i])[0]     #tidx1600[i]=ut.find_predecessor(allmaps['aia1600']['time1600'],vla0['vla0']['timevla'][i])[0]     #tidx335[i]=ut.find_predecessor(allmaps['aia335']['time335'],vla0['vla0']['timevla'][i])[0]     #tidx171[i]=ut.find_predecessor(allmaps['aia171']['time171'],vla0['vla0']['timevla'][i])[0]     #tidx131[i]=ut.find_predecessor(allmaps['aia131']['time131'],vla0['vla0']['timevla'][i])[0]     #tidx94[i]=ut.find_predecessor(allmaps['aia94']['time94'],vla0['vla0']['timevla'][i])[0]     tidx1700[i]=ut.find_predecessor(allmaps['aia1700']['time1700'],timevla_all1[i])[0]     tidx1600[i]=ut.find_predecessor(allmaps['aia1600']['time1600'],timevla_all1[i])[0]     tidx335[i]=ut.find_predecessor(allmaps['aia335']['time335'],timevla_all1[i])[0]     tidx171[i]=ut.find_predecessor(allmaps['aia171']['time171'],timevla_all1[i])[0]     tidx131[i]=ut.find_predecessor(allmaps['aia131']['time131'],timevla_all1[i])[0]     tidx94[i]=ut.find_predecessor(allmaps['aia94']['time94'],timevla_all1[i])[0] for i in range(m): tidx335=[0]*m;tidx1600=[0]*m;tidx1700=[0]*m tidx94=[0]*m;tidx131=[0]*m;tidx171=[0]*m m=len(timevla_all1) Tb_mean_r1=Tb0[:,:,115:145,115:145].mean(axis=(2,3)) #Tb_mean_r1=Tb[:,:,30:80,115:145].mean(axis=(2,3)) Tbmax_ds=Tb0.max(axis=(2,3)) Tb7=np.array(vla7['vla7']['datavla']).reshape(1,2399,256,256) #Tb6=np.array(vla6['vla6']['datavla']).reshape(1,2399,256,256) #Tb5=np.array(vla5['vla5']['datavla']).reshape(1,2399,256,256) #Tb4=np.array(vla4['vla4']['datavla']).reshape(1,2399,256,256) #Tb3=np.array(vla3['vla3']['datavla']).reshape(1,2399,256,256) #Tb2=np.array(vla2['vla2']['datavla']).reshape(1,2399,256,256) #Tb1=np.array(vla1['vla1']['datavla']).reshape(1,2399,256,256) Tb0=np.array(vla0['vla0']['datavla']).reshape(1,2399,256,256) #Tb=np.array(allmaps['vla']['datavla']).reshape(32,119,150,200) ################# Analysis ################# freq=np.linspace(0.997,1.245,32) timed1600=allmaps['aiad1600']['timed1600'];timed1700=allmaps['aiad1700']['timed1700'];time171=allmaps['aiad171']['timed171'] timed94=allmaps['aiad94']['timed94'];timed131=allmaps['aiad131']['timed131'];time335=allmaps['aiad335']['timed335'] time1600=allmaps['aia1600']['time1600'];time1700=allmaps['aia1700']['time1700'];time171=allmaps['aia171']['time171'] time94=allmaps['aia94']['time94'];time131=allmaps['aia131']['time131'];time335=allmaps['aia335']['time335'] timevla=vla0['vla0']['timevla']  #vla7=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_7_50ms.p','rb')) #vla6=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_6_50ms.p','rb')) #vla5=pickle.load(open('/medi8a/rohit/VLA/20160409/20160409_vla_spw_5_50ms.p','rb')) #vla4=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_4_50ms.p','rb')) print "Reading 5 and 7.." #vla3=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_3_50ms.p','rb')) #vla2=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_2_50ms.p','rb')) #vla1=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_1_50ms.p','rb')) vla0=pickle.load(open('/media/rohit/VLA/20160409/20160409_vla_spw_0_50ms.p','rb')) allmaps=pickle.load(open('/media/rohit/VLA/20160409/20160409_submap_aia_50ms.p','rb')) ################ Read submaps ##############            timstr_171[i]= list171[i].split('T')[-1].split('Z')[0] ad     �     e       �  �  a  )  �  �  z  V  /  .  -  �  �  �  �  �  �  <  �  �  �  �  �  �  a  B  .         �  �  �  �  e  =  1    �
  �
  �
  q
  p
  B
  A
  �	  �	  d	  	  �  n    �  �  �  �  9  �  �  �  �  �  Y  A  $          �  �  -    �  �  �  s  a  P  G  4  #    �  �  t  s  c  7    �  �  *  )  (  '    �  �  �  �  �                            if(plot_euv_time): plot_euv_time=1  ################ PLOTTING ################### sys.exit()    ds_LL1=np.hstack((ds1s,np.subtract(ds1s[:,-1],-1*ds_LL[6:512].swapaxes(0,1)+28).swapaxes(0,1))) ds1s=np.subtract(ds1['spec'][0][0].swapaxes(0,1),ds1['spec'][0][0][:,0]).swapaxes(0,1)/3  freq=freq.swapaxes(0,1).flatten()/1.e9 ds_RR=ds[1].swapaxes(0,1).reshape(512,2400) ds_LL=ds[0].swapaxes(0,1).reshape(512,2400) ds=np.array(ds)              ds[i][j][k]=np.hstack((ds_[i,j,2089*k:2089*(k+1)],ds_[i,j,16712+k*311:16712+(k+1)*311]))         for k in range(8):         ds[i][j]=[0]*8     for j in range(64):     ds[i]=[0]*64 for i in range(2): ds=[0]*2 ds_=ds_[:,0,:,:] tim=np.array(tim)     tim[i]=np.hstack((tim_[2089*i:2089*(i+1)],tim_[16712+i*311:16712+(i+1)*311])) for i in range(8): tim=[0]*8 tim_=data['tim'];freq=data['freq'];ds_=data['spec'] data=np.load(specfile) specfile='/media/rohit/VLA/20160409/sun_L_20160409T1844-1846UT.50ms.cal.ms.dspec.median.npz' ds1=np.load('/media/rohit/VLA/20160409/sun_L_20160409T184000-184400UT.50ms.cal.ms.dspec.npz') ############### MAKE DS #####################    plt.show() plt.plot(fmtime,fmrate,'o-') fmtime=fmtime-fmtime[0] fmrate=fm1.data['RATE'];fmtime=fm1.data['TIME'] fm0=fm[0];fm1=fm[1] fm=fits.open('/home/i4ds1807205/Dropbox/20160409/fermi/glg_cspec_n5_160409_v00_data.fits')   gf0540=goes['lx'][1];gf1080=goes['lx'][0];gtime=goes['tarray'] goes=readsav('/home/i4ds1807205/Dropbox/20160409/fermi/idlsave_goes.sav') ################ FERMI & GOES & VLA DS #######################       tidx1700[i]=ut.find_predecessor(allmaps['aia1700']['time1700'],timevla[i][0])[0]     tidx1600[i]=ut.find_predecessor(allmaps['aia1600']['time1600'],timevla[i][0])[0]     tidx335[i]=ut.find_predecessor(allmaps['aia335']['time335'],timevla[i][0])[0]     tidx171[i]=ut.find_predecessor(allmaps['aia171']['time171'],timevla[i][0])[0]     tidx131[i]=ut.find_predecessor(allmaps['aia131']['time131'],timevla[i][0])[0]     tidx94[i]=ut.find_predecessor(allmaps['aia94']['time94'],timevla[i][0])[0] for i in range(2000): tidx94=[0]*2000;tidx131=[0]*2000;tidx171=[0]*2000;tidx193=[0]*2000;tidx335=[0]*2000;tidx1600=[0]*2000;tidx1700=[0]*2000  #############################################  ts1700=get_ts(data1700,350,500,600,750) ts1600=get_ts(data1600,350,500,600,750) ts335=get_ts(data335,350,500,600,750) ts131=get_ts(data131,350,500,600,750) ts94=get_ts(data94,350,500,600,750) #Timeseries data1700=allmaps['aia1700']['data1700'] data1600=allmaps['aia1600']['data1600'] data335=allmaps['aia335']['data335'] data171=allmaps['aia171']['data171'] data131=allmaps['aia131']['data131'] data94=allmaps['aia94']['data94']       return ts     ts=np.array(ts)         ts[i]=np.nanmean(d[i])         #ts[i]=np.nanmax(d[i][xl:xr,yl:yr])     for i in range(len(d)):     ts=[0]*len(d) def get_ts(d,xl,xr,yl,yr):  Tb_r=np.array(Tb_r)         Tb_r[i][j]=np.mean(datavla_v[j][0][re[i][0]:re[i][1],re[i][2]:re[i][3]])         #Tb_r[i][j]=np.mean(Tb1[0][j][re[i][0]:re[i][1],re[i][2]:re[i][3]])     for j in range(2000):     Tb_r[i]=[0]*2000 for i in range(5): Tb_r=[0]*5  re=[[124,134,120,130],[140,150,90,100],[95,115,70,90],[105,125,30,50],[95,115,95,115]]   vlasize_fwhm[np.isnan(vlasize_fwhm)]=0 vlasize_fwhm=np.array(vlasize_fwhm) vlasize=np.array(vlasize)             vlasize_fwhm[k][i][j]=bimage_fwhm[np.isfinite(bimage_fwhm)].sum()*2.0             vlasize[k][i][j]=bimage[np.isfinite(bimage)].sum()*2.0             bimage_fwhm=ut.get_bimage(Tb0[i][j],lev[k])             bimage=ut.get_bimage(Tb0[i][j],lev[k]*3.e7/np.nanmax(Tb0[i][j]))         for j in range(Tb0.shape[1]):         vlasize_fwhm[k][i]=[0]*Tb0.shape[1] ad  s  7     *       (  �  �  d  $  �  �  �  y  .  �  �  w  '  �
  �
  �
  �
  �
  �
  i
  8
  �	  �	  �	  �	  �	  w	  U	  }  :  �  �      �  y  �  �    �  7  �  �  �  �  �  X  	  �  �  q    �  �  Y  (  �  �  m  B  A                                                        ax[2].set_xlabel('Time (HH:MM:SS UT)')     ax[2].set_xticks([0,30,60,90,120]);ax[2].set_xticklabels(['18:44:00','18:44:30','18:45:00','18:45:30','18:46:00'])     ax[2].legend()     ax[2].plot(vlasize[3,10],'o-',label='27 MK')     ax[2].plot(vlasize[2,10],'o-',label='21 MK')     #ax[2].plot(vlasize[1,10],'o-',label='18 MK')     ax[2].plot(vlasize[0,10],'o-',label='15 MK (1.ax0.text(xlaia+10,ylaia+10,str(np.round(v6.meta['restfrq']/1.e9,3))+' MHz',fontsize=12,color=color_array[0][0:aaaaaaaaaaaaax0.text(-900+10,100+10,str(np.round(v6.meta['restfrq']/1.e9,3))+' GHz',fontsize=18,color=color_array[50][0:3]) ax0.text(-900+10,100+20,str(np.round(v4.meta['restfrq']/1.e9,3))+' GHz',fontsize=18,color=color_array[40][0:3]) ax0.text(-900+10,100+30,str(np.round(v2.meta['restfrq']/1.e9,3))+' GHz',fontsize=18,color=color_array[30][0:3]) ax0.text(-900+10,100+40,str(np.round(dd.meta['restfrq']/1.e9,3))+' GHz',fontsize=18,color=color_array[0][0:3]) v6.draw_contours(levels=lev1,colors=color_array[50][0:3],linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) v4.draw_contours(levels=lev1,colors=color_array[40][0:3],linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) v2.draw_contours(levels=lev1,colors=color_array[30][0:3],linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) dd.draw_contours(levels=lev1,colors=color_array[0][0:3],linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2) lev1=np.array([70,75,85,95])*u.percent #lev1=(1.5e7/dd.data.max())*np.array([60,70,80,90])*u.percent p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2) dd=v;dd.data[np.isnan(dd.data)]=0 cc=maphmi[-1] ax0 = f.add_subplot(111) f=plt.figure(figsize=(10,10))  plt.register_cmap(cmap=map_object) map_object = LinearSegmentedColormap.from_list(name='rainbow_alpha',colors=color_array) color_array[:,-1] = np.linspace(0.0,1.0,ncolors) color_array = plt.get_cmap('gist_rainbow')(range(ncolors)) ncolors = 256 from matplotlib.colors import LinearSegmentedColormap   plt.show() ax0.set_xlim([-900,-700]),ax0.set_ylim([100,300]) #ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow') #ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r') #ax0.plot(b_hp_fr.Tx,b_hp_fr.Ty,'o',markersize=3) #ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia]) ax0.set_title('AIA 171 $\AA$:18:42:10 UT VLA: 18:44:43.00-18:44:43.05 UT') dd.draw_contours(levels=lev1,colors='r',linewidths=2,extent=[xlvla,xrvla,ylvla,yrvla])#[xlpix,xrpix,ylpix,yrpix]) xlvla=dd.center.Tx.value-2.0*int(dd.data.shape[0]/2);xrvla=dd.center.Tx.value+2.0*int(dd.data.shape[0]/2);ylvla=dd.center.Ty.value-2.0*int(dd.data.shape[1]/2);yrvla=dd.center.Ty.value+2.0*int(dd.data.shape[0]/2) lev1=np.array([60,70,80,90])*u.percent #lev1=(1.5e7/dd.data.max())*np.array([60,70,80,90])*u.percent ax0.plot(b_hp_ls[0],b_hp_ls[1],'o',markersize=2,color='orange') ax0.plot(b_hp_fr[0],b_hp_fr[1],'o',markersize=2,color='magenta') ax0.plot(b_hp_euv[0],b_hp_euv[1],'o',markersize=2,color='cyan') p=cc.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto') xlaia=cc.center.Tx.value-0.61*int(cc.data.shape[0]/2);xraia=cc.center.Tx.value+0.61*int(cc.data.shape[0]/2);ylaia=cc.center.Ty.value-0.61*int(cc.data.shape[1]/2);yraia=cc.center.Ty.value+0.61*int(cc.data.shape[0]/2) ad  /
  �
            �  |  ,  �  �  b             �  �  z  Q    �  �  9  �  �  �  h  U  �
  �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ax[2].set_xlabel('Time (HH:MM:SS UT)')     ax[2].set_xticks([0,30,60,90,120]);ax[2].set_xticklabels(['18:44:00','18:44:30','18:45:00','18:45:30','18:46:00'])     ax[2].legend()     ax[2].plot(vlasize[3,10],'o-',label='27 MK')     ax[2].plot(vlasize[2,10],'o-',label='21 MK')     #ax[2].plot(vlasize[1,10],'o-',label='18 MK')     ax[2].plot(vlasize[0,10],'o-',label='15 MK (1.077 GHz)')     ax[1].plot(Tb_mean_r1[10]/1.e6,'o-',label='1.077 GHz');ax[1].legend()     ax[0].set_yticks([0,10,20,30]);ax[0].set_yticklabels([freq[0],freq[10],freq[20],freq[30]])     fig.colorbar(im0,cax=cax,label='T$_{B}$ (MK)')     cax = divider.append_axes('right', size='5%', pad=0.05)     divider = make_axes_locatable(ax[0])     im0=ax[0].imshow(Tb_mean_r1/1.e6,origin=0,cmap='jet',interpolation='None')     fig,ax=plt.subplots(3,1,sharex=True) if(plot_vlasize): plot_vlasize=1   plt.show() ax0.set_title('HMI: 18:50:47 UT VLA: 18:44:43.00-18:44:43.05 UT') p=ee.plot(axes=ax0,extent=[xlaia,xraia,ylaia,yraia],aspect='auto',cmap='rainbow_alpha',vmin=100,vmax=8000,alpha=0.7) ee=allmaps['aia171']['map171'][10] ax0.set_xlim([-900,-700]),ax0.set_ylim([100,300]) #ax0.text(-1200,50,'Contours: 3, 4.5, 6, 7.5, 9, 10, 12, 13 MK',color='yellow') #ax0.text(-1200,0,str(np.round(dd.meta['crval3']/1.e9,4))+' GHz',color='r') ax0.set_xlim([xlaia,xraia]);ax0.set_ylim([ylaia,yraia]) 